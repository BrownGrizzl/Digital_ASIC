module add_signed_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [22:0] A;
  input [12:0] B;
  output [23:0] Z;
  wire [22:0] A;
  wire [12:0] B;
  wire [23:0] Z;
  wire n_66, n_67, n_68, n_69, n_70, n_73, n_74, n_75;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  not g3 (Z[23], n_73);
  nand g4 (n_75, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_66, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_67, A[9], B[9]);
  nand g59 (n_68, A[9], n_66);
  nand g60 (n_69, B[9], n_66);
  nand g61 (n_119, n_67, n_68, n_69);
  xor g62 (n_70, A[9], B[9]);
  xor g63 (Z[9], n_66, n_70);
  nand g64 (n_74, A[10], B[10]);
  nand g65 (n_120, A[10], n_119);
  nand g66 (n_121, B[10], n_119);
  nand g67 (n_123, n_74, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_119, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[12]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[12], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[12]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[12]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[12], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[12]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[12]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[12], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[12]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[12]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[12], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[12]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[12]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[12], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[12]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[12]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[12], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[12]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[19], B[12]);
  nand g119 (n_165, A[19], n_163);
  nand g120 (n_166, B[12], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[19], B[12]);
  xor g123 (Z[19], n_163, n_167);
  nand g124 (n_169, A[20], B[12]);
  nand g125 (n_170, A[20], n_168);
  nand g126 (n_171, B[12], n_168);
  nand g127 (n_173, n_169, n_170, n_171);
  xor g128 (n_172, A[20], B[12]);
  xor g129 (Z[20], n_168, n_172);
  nand g130 (n_174, A[21], B[12]);
  nand g131 (n_175, A[21], n_173);
  nand g132 (n_176, B[12], n_173);
  nand g133 (n_178, n_174, n_175, n_176);
  xor g134 (n_177, A[21], B[12]);
  xor g135 (Z[21], n_173, n_177);
  nand g139 (n_73, n_179, n_180, n_181);
  xor g141 (Z[22], n_178, n_182);
  or g143 (n_179, A[22], B[12]);
  xor g144 (n_182, A[22], B[12]);
  or g145 (n_81, wc, n_75);
  not gc (wc, A[1]);
  or g146 (n_82, wc0, n_75);
  not gc0 (wc0, B[1]);
  xnor g147 (Z[1], n_75, n_83);
  or g148 (n_180, A[22], wc1);
  not gc1 (wc1, n_178);
  or g149 (n_181, B[12], wc2);
  not gc2 (wc2, n_178);
endmodule

module add_signed_GENERIC(A, B, Z);
  input [22:0] A;
  input [12:0] B;
  output [23:0] Z;
  wire [22:0] A;
  wire [12:0] B;
  wire [23:0] Z;
  add_signed_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_23_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [15:0] A;
  input [16:0] B;
  output [16:0] Z;
  wire [15:0] A;
  wire [16:0] B;
  wire [16:0] Z;
  wire n_54, n_57, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_139;
  nand g4 (n_57, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_62, A[1], B[1]);
  nand g13 (n_66, n_62, n_63, n_64);
  xor g14 (n_65, A[1], B[1]);
  nand g16 (n_67, A[2], B[2]);
  nand g17 (n_68, A[2], n_66);
  nand g18 (n_69, B[2], n_66);
  nand g19 (n_71, n_67, n_68, n_69);
  xor g20 (n_70, A[2], B[2]);
  xor g21 (Z[2], n_66, n_70);
  nand g22 (n_72, A[3], B[3]);
  nand g23 (n_73, A[3], n_71);
  nand g24 (n_74, B[3], n_71);
  nand g25 (n_76, n_72, n_73, n_74);
  xor g26 (n_75, A[3], B[3]);
  xor g27 (Z[3], n_71, n_75);
  nand g28 (n_77, A[4], B[4]);
  nand g29 (n_78, A[4], n_76);
  nand g30 (n_79, B[4], n_76);
  nand g31 (n_81, n_77, n_78, n_79);
  xor g32 (n_80, A[4], B[4]);
  xor g33 (Z[4], n_76, n_80);
  nand g34 (n_82, A[5], B[5]);
  nand g35 (n_83, A[5], n_81);
  nand g36 (n_84, B[5], n_81);
  nand g37 (n_86, n_82, n_83, n_84);
  xor g38 (n_85, A[5], B[5]);
  xor g39 (Z[5], n_81, n_85);
  nand g40 (n_87, A[6], B[6]);
  nand g41 (n_88, A[6], n_86);
  nand g42 (n_89, B[6], n_86);
  nand g43 (n_91, n_87, n_88, n_89);
  xor g44 (n_90, A[6], B[6]);
  xor g45 (Z[6], n_86, n_90);
  nand g46 (n_92, A[7], B[7]);
  nand g47 (n_54, A[7], n_91);
  nand g48 (n_93, B[7], n_91);
  nand g49 (n_95, n_92, n_54, n_93);
  xor g50 (n_94, A[7], B[7]);
  xor g51 (Z[7], n_91, n_94);
  nand g52 (n_96, A[8], B[8]);
  nand g53 (n_97, A[8], n_95);
  nand g54 (n_98, B[8], n_95);
  nand g55 (n_100, n_96, n_97, n_98);
  xor g56 (n_99, A[8], B[8]);
  xor g57 (Z[8], n_95, n_99);
  nand g58 (n_101, A[9], B[9]);
  nand g59 (n_102, A[9], n_100);
  nand g60 (n_103, B[9], n_100);
  nand g61 (n_105, n_101, n_102, n_103);
  xor g62 (n_104, A[9], B[9]);
  xor g63 (Z[9], n_100, n_104);
  nand g64 (n_106, A[10], B[10]);
  nand g65 (n_107, A[10], n_105);
  nand g66 (n_108, B[10], n_105);
  nand g67 (n_110, n_106, n_107, n_108);
  xor g68 (n_109, A[10], B[10]);
  xor g69 (Z[10], n_105, n_109);
  nand g70 (n_111, A[11], B[11]);
  nand g71 (n_112, A[11], n_110);
  nand g72 (n_113, B[11], n_110);
  nand g73 (n_115, n_111, n_112, n_113);
  xor g74 (n_114, A[11], B[11]);
  xor g75 (Z[11], n_110, n_114);
  nand g76 (n_116, A[12], B[12]);
  nand g77 (n_117, A[12], n_115);
  nand g78 (n_118, B[12], n_115);
  nand g79 (n_120, n_116, n_117, n_118);
  xor g80 (n_119, A[12], B[12]);
  xor g81 (Z[12], n_115, n_119);
  nand g82 (n_121, A[13], B[13]);
  nand g83 (n_122, A[13], n_120);
  nand g84 (n_123, B[13], n_120);
  nand g85 (n_125, n_121, n_122, n_123);
  xor g86 (n_124, A[13], B[13]);
  xor g87 (Z[13], n_120, n_124);
  nand g88 (n_126, A[14], B[14]);
  nand g89 (n_127, A[14], n_125);
  nand g90 (n_128, B[14], n_125);
  nand g91 (n_130, n_126, n_127, n_128);
  xor g92 (n_129, A[14], B[14]);
  xor g93 (Z[14], n_125, n_129);
  nand g94 (n_131, A[15], B[15]);
  nand g95 (n_132, A[15], n_130);
  nand g96 (n_133, B[15], n_130);
  nand g97 (n_135, n_131, n_132, n_133);
  xor g98 (n_134, A[15], B[15]);
  xor g99 (Z[15], n_130, n_134);
  xor g105 (Z[16], n_135, n_139);
  xor g107 (n_139, A[15], B[16]);
  or g108 (n_63, wc, n_57);
  not gc (wc, A[1]);
  or g109 (n_64, wc0, n_57);
  not gc0 (wc0, B[1]);
  xnor g110 (Z[1], n_57, n_65);
endmodule

module add_signed_23_GENERIC(A, B, Z);
  input [15:0] A;
  input [16:0] B;
  output [16:0] Z;
  wire [15:0] A;
  wire [16:0] B;
  wire [16:0] Z;
  add_signed_23_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_24_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [18:0] A;
  input [21:0] B;
  output [21:0] Z;
  wire [18:0] A;
  wire [21:0] B;
  wire [21:0] Z;
  wire n_67, n_68, n_69, n_72, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_177;
  nand g4 (n_72, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_67, A[9], B[9]);
  nand g59 (n_68, A[9], n_116);
  nand g60 (n_69, B[9], n_116);
  nand g61 (n_118, n_67, n_68, n_69);
  xor g62 (n_117, A[9], B[9]);
  xor g63 (Z[9], n_116, n_117);
  nand g64 (n_119, A[10], B[10]);
  nand g65 (n_120, A[10], n_118);
  nand g66 (n_121, B[10], n_118);
  nand g67 (n_123, n_119, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_118, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[13]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[13], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[13]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[14]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[14], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[14]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[15]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[15], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[15]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[16]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[16], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[16]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[17]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[17], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[17]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[18]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[18], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[18]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[18], B[19]);
  nand g119 (n_165, A[18], n_163);
  nand g120 (n_166, B[19], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[18], B[19]);
  xor g123 (Z[19], n_163, n_167);
  nand g124 (n_169, A[18], B[20]);
  nand g125 (n_170, A[18], n_168);
  nand g126 (n_171, B[20], n_168);
  nand g127 (n_173, n_169, n_170, n_171);
  xor g128 (n_172, A[18], B[20]);
  xor g129 (Z[20], n_168, n_172);
  xor g135 (Z[21], n_173, n_177);
  xor g137 (n_177, A[18], B[21]);
  or g138 (n_78, wc, n_72);
  not gc (wc, A[1]);
  or g139 (n_79, wc0, n_72);
  not gc0 (wc0, B[1]);
  xnor g140 (Z[1], n_72, n_80);
endmodule

module add_signed_24_GENERIC(A, B, Z);
  input [18:0] A;
  input [21:0] B;
  output [21:0] Z;
  wire [18:0] A;
  wire [21:0] B;
  wire [21:0] Z;
  add_signed_24_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_25_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [22:0] A;
  input [18:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [18:0] B;
  wire [22:0] Z;
  wire n_69, n_70, n_75, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_186;
  nand g4 (n_75, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_69, B[9], n_119);
  nand g61 (n_122, n_120, n_121, n_69);
  xor g62 (n_70, A[9], B[9]);
  xor g63 (Z[9], n_119, n_70);
  nand g64 (n_123, A[10], B[10]);
  nand g65 (n_124, A[10], n_122);
  nand g66 (n_125, B[10], n_122);
  nand g67 (n_127, n_123, n_124, n_125);
  xor g68 (n_126, A[10], B[10]);
  xor g69 (Z[10], n_122, n_126);
  nand g70 (n_128, A[11], B[11]);
  nand g71 (n_129, A[11], n_127);
  nand g72 (n_130, B[11], n_127);
  nand g73 (n_132, n_128, n_129, n_130);
  xor g74 (n_131, A[11], B[11]);
  xor g75 (Z[11], n_127, n_131);
  nand g76 (n_133, A[12], B[12]);
  nand g77 (n_134, A[12], n_132);
  nand g78 (n_135, B[12], n_132);
  nand g79 (n_137, n_133, n_134, n_135);
  xor g80 (n_136, A[12], B[12]);
  xor g81 (Z[12], n_132, n_136);
  nand g82 (n_138, A[13], B[13]);
  nand g83 (n_139, A[13], n_137);
  nand g84 (n_140, B[13], n_137);
  nand g85 (n_142, n_138, n_139, n_140);
  xor g86 (n_141, A[13], B[13]);
  xor g87 (Z[13], n_137, n_141);
  nand g88 (n_143, A[14], B[14]);
  nand g89 (n_144, A[14], n_142);
  nand g90 (n_145, B[14], n_142);
  nand g91 (n_147, n_143, n_144, n_145);
  xor g92 (n_146, A[14], B[14]);
  xor g93 (Z[14], n_142, n_146);
  nand g94 (n_148, A[15], B[15]);
  nand g95 (n_149, A[15], n_147);
  nand g96 (n_150, B[15], n_147);
  nand g97 (n_152, n_148, n_149, n_150);
  xor g98 (n_151, A[15], B[15]);
  xor g99 (Z[15], n_147, n_151);
  nand g100 (n_153, A[16], B[16]);
  nand g101 (n_154, A[16], n_152);
  nand g102 (n_155, B[16], n_152);
  nand g103 (n_157, n_153, n_154, n_155);
  xor g104 (n_156, A[16], B[16]);
  xor g105 (Z[16], n_152, n_156);
  nand g106 (n_158, A[17], B[17]);
  nand g107 (n_159, A[17], n_157);
  nand g108 (n_160, B[17], n_157);
  nand g109 (n_162, n_158, n_159, n_160);
  xor g110 (n_161, A[17], B[17]);
  xor g111 (Z[17], n_157, n_161);
  nand g112 (n_163, A[18], B[18]);
  nand g113 (n_164, A[18], n_162);
  nand g114 (n_165, B[18], n_162);
  nand g115 (n_167, n_163, n_164, n_165);
  xor g116 (n_166, A[18], B[18]);
  xor g117 (Z[18], n_162, n_166);
  nand g118 (n_168, A[19], B[18]);
  nand g119 (n_169, A[19], n_167);
  nand g120 (n_170, B[18], n_167);
  nand g121 (n_172, n_168, n_169, n_170);
  xor g122 (n_171, A[19], B[18]);
  xor g123 (Z[19], n_167, n_171);
  nand g124 (n_173, A[20], B[18]);
  nand g125 (n_174, A[20], n_172);
  nand g126 (n_175, B[18], n_172);
  nand g127 (n_177, n_173, n_174, n_175);
  xor g128 (n_176, A[20], B[18]);
  xor g129 (Z[20], n_172, n_176);
  nand g130 (n_178, A[21], B[18]);
  nand g131 (n_179, A[21], n_177);
  nand g132 (n_180, B[18], n_177);
  nand g133 (n_182, n_178, n_179, n_180);
  xor g134 (n_181, A[21], B[18]);
  xor g135 (Z[21], n_177, n_181);
  xor g141 (Z[22], n_182, n_186);
  xor g143 (n_186, A[22], B[18]);
  or g144 (n_81, wc, n_75);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_75);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_75, n_83);
endmodule

module add_signed_25_GENERIC(A, B, Z);
  input [22:0] A;
  input [18:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [18:0] B;
  wire [22:0] Z;
  add_signed_25_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_26_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [22:0] A;
  input [14:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [14:0] B;
  wire [22:0] Z;
  wire n_66, n_67, n_68, n_69, n_70, n_75, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_183;
  nand g4 (n_75, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_66, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_67, A[9], B[9]);
  nand g59 (n_68, A[9], n_66);
  nand g60 (n_69, B[9], n_66);
  nand g61 (n_119, n_67, n_68, n_69);
  xor g62 (n_70, A[9], B[9]);
  xor g63 (Z[9], n_66, n_70);
  nand g64 (n_120, A[10], B[10]);
  nand g65 (n_121, A[10], n_119);
  nand g66 (n_122, B[10], n_119);
  nand g67 (n_124, n_120, n_121, n_122);
  xor g68 (n_123, A[10], B[10]);
  xor g69 (Z[10], n_119, n_123);
  nand g70 (n_125, A[11], B[11]);
  nand g71 (n_126, A[11], n_124);
  nand g72 (n_127, B[11], n_124);
  nand g73 (n_129, n_125, n_126, n_127);
  xor g74 (n_128, A[11], B[11]);
  xor g75 (Z[11], n_124, n_128);
  nand g76 (n_130, A[12], B[12]);
  nand g77 (n_131, A[12], n_129);
  nand g78 (n_132, B[12], n_129);
  nand g79 (n_134, n_130, n_131, n_132);
  xor g80 (n_133, A[12], B[12]);
  xor g81 (Z[12], n_129, n_133);
  nand g82 (n_135, A[13], B[13]);
  nand g83 (n_136, A[13], n_134);
  nand g84 (n_137, B[13], n_134);
  nand g85 (n_139, n_135, n_136, n_137);
  xor g86 (n_138, A[13], B[13]);
  xor g87 (Z[13], n_134, n_138);
  nand g88 (n_140, A[14], B[14]);
  nand g89 (n_141, A[14], n_139);
  nand g90 (n_142, B[14], n_139);
  nand g91 (n_144, n_140, n_141, n_142);
  xor g92 (n_143, A[14], B[14]);
  xor g93 (Z[14], n_139, n_143);
  nand g94 (n_145, A[15], B[14]);
  nand g95 (n_146, A[15], n_144);
  nand g96 (n_147, B[14], n_144);
  nand g97 (n_149, n_145, n_146, n_147);
  xor g98 (n_148, A[15], B[14]);
  xor g99 (Z[15], n_144, n_148);
  nand g100 (n_150, A[16], B[14]);
  nand g101 (n_151, A[16], n_149);
  nand g102 (n_152, B[14], n_149);
  nand g103 (n_154, n_150, n_151, n_152);
  xor g104 (n_153, A[16], B[14]);
  xor g105 (Z[16], n_149, n_153);
  nand g106 (n_155, A[17], B[14]);
  nand g107 (n_156, A[17], n_154);
  nand g108 (n_157, B[14], n_154);
  nand g109 (n_159, n_155, n_156, n_157);
  xor g110 (n_158, A[17], B[14]);
  xor g111 (Z[17], n_154, n_158);
  nand g112 (n_160, A[18], B[14]);
  nand g113 (n_161, A[18], n_159);
  nand g114 (n_162, B[14], n_159);
  nand g115 (n_164, n_160, n_161, n_162);
  xor g116 (n_163, A[18], B[14]);
  xor g117 (Z[18], n_159, n_163);
  nand g118 (n_165, A[19], B[14]);
  nand g119 (n_166, A[19], n_164);
  nand g120 (n_167, B[14], n_164);
  nand g121 (n_169, n_165, n_166, n_167);
  xor g122 (n_168, A[19], B[14]);
  xor g123 (Z[19], n_164, n_168);
  nand g124 (n_170, A[20], B[14]);
  nand g125 (n_171, A[20], n_169);
  nand g126 (n_172, B[14], n_169);
  nand g127 (n_174, n_170, n_171, n_172);
  xor g128 (n_173, A[20], B[14]);
  xor g129 (Z[20], n_169, n_173);
  nand g130 (n_175, A[21], B[14]);
  nand g131 (n_176, A[21], n_174);
  nand g132 (n_177, B[14], n_174);
  nand g133 (n_179, n_175, n_176, n_177);
  xor g134 (n_178, A[21], B[14]);
  xor g135 (Z[21], n_174, n_178);
  xor g141 (Z[22], n_179, n_183);
  xor g143 (n_183, A[22], B[14]);
  or g144 (n_81, wc, n_75);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_75);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_75, n_83);
endmodule

module add_signed_26_GENERIC(A, B, Z);
  input [22:0] A;
  input [14:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [14:0] B;
  wire [22:0] Z;
  add_signed_26_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_303_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  wire n_71, n_72, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180;
  not g3 (Z[22], n_71);
  nand g4 (n_72, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  nand g133 (n_71, n_177, n_178, n_179);
  xor g135 (Z[21], n_176, n_180);
  or g137 (n_177, A[21], B[21]);
  xor g138 (n_180, A[21], B[21]);
  or g139 (n_78, wc, n_72);
  not gc (wc, A[1]);
  or g140 (n_79, wc0, n_72);
  not gc0 (wc0, B[1]);
  xnor g141 (Z[1], n_72, n_80);
  or g142 (n_178, A[21], wc1);
  not gc1 (wc1, n_176);
  or g143 (n_179, B[21], wc2);
  not gc2 (wc2, n_176);
endmodule

module add_signed_303_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  add_signed_303_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_6_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [22:0] A;
  input [16:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [16:0] B;
  wire [22:0] Z;
  wire n_67, n_68, n_69, n_70, n_75, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_184;
  nand g4 (n_75, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_67, A[9], B[9]);
  nand g59 (n_68, A[9], n_119);
  nand g60 (n_69, B[9], n_119);
  nand g61 (n_120, n_67, n_68, n_69);
  xor g62 (n_70, A[9], B[9]);
  xor g63 (Z[9], n_119, n_70);
  nand g64 (n_121, A[10], B[10]);
  nand g65 (n_122, A[10], n_120);
  nand g66 (n_123, B[10], n_120);
  nand g67 (n_125, n_121, n_122, n_123);
  xor g68 (n_124, A[10], B[10]);
  xor g69 (Z[10], n_120, n_124);
  nand g70 (n_126, A[11], B[11]);
  nand g71 (n_127, A[11], n_125);
  nand g72 (n_128, B[11], n_125);
  nand g73 (n_130, n_126, n_127, n_128);
  xor g74 (n_129, A[11], B[11]);
  xor g75 (Z[11], n_125, n_129);
  nand g76 (n_131, A[12], B[12]);
  nand g77 (n_132, A[12], n_130);
  nand g78 (n_133, B[12], n_130);
  nand g79 (n_135, n_131, n_132, n_133);
  xor g80 (n_134, A[12], B[12]);
  xor g81 (Z[12], n_130, n_134);
  nand g82 (n_136, A[13], B[13]);
  nand g83 (n_137, A[13], n_135);
  nand g84 (n_138, B[13], n_135);
  nand g85 (n_140, n_136, n_137, n_138);
  xor g86 (n_139, A[13], B[13]);
  xor g87 (Z[13], n_135, n_139);
  nand g88 (n_141, A[14], B[14]);
  nand g89 (n_142, A[14], n_140);
  nand g90 (n_143, B[14], n_140);
  nand g91 (n_145, n_141, n_142, n_143);
  xor g92 (n_144, A[14], B[14]);
  xor g93 (Z[14], n_140, n_144);
  nand g94 (n_146, A[15], B[15]);
  nand g95 (n_147, A[15], n_145);
  nand g96 (n_148, B[15], n_145);
  nand g97 (n_150, n_146, n_147, n_148);
  xor g98 (n_149, A[15], B[15]);
  xor g99 (Z[15], n_145, n_149);
  nand g100 (n_151, A[16], B[16]);
  nand g101 (n_152, A[16], n_150);
  nand g102 (n_153, B[16], n_150);
  nand g103 (n_155, n_151, n_152, n_153);
  xor g104 (n_154, A[16], B[16]);
  xor g105 (Z[16], n_150, n_154);
  nand g106 (n_156, A[17], B[16]);
  nand g107 (n_157, A[17], n_155);
  nand g108 (n_158, B[16], n_155);
  nand g109 (n_160, n_156, n_157, n_158);
  xor g110 (n_159, A[17], B[16]);
  xor g111 (Z[17], n_155, n_159);
  nand g112 (n_161, A[18], B[16]);
  nand g113 (n_162, A[18], n_160);
  nand g114 (n_163, B[16], n_160);
  nand g115 (n_165, n_161, n_162, n_163);
  xor g116 (n_164, A[18], B[16]);
  xor g117 (Z[18], n_160, n_164);
  nand g118 (n_166, A[19], B[16]);
  nand g119 (n_167, A[19], n_165);
  nand g120 (n_168, B[16], n_165);
  nand g121 (n_170, n_166, n_167, n_168);
  xor g122 (n_169, A[19], B[16]);
  xor g123 (Z[19], n_165, n_169);
  nand g124 (n_171, A[20], B[16]);
  nand g125 (n_172, A[20], n_170);
  nand g126 (n_173, B[16], n_170);
  nand g127 (n_175, n_171, n_172, n_173);
  xor g128 (n_174, A[20], B[16]);
  xor g129 (Z[20], n_170, n_174);
  nand g130 (n_176, A[21], B[16]);
  nand g131 (n_177, A[21], n_175);
  nand g132 (n_178, B[16], n_175);
  nand g133 (n_180, n_176, n_177, n_178);
  xor g134 (n_179, A[21], B[16]);
  xor g135 (Z[21], n_175, n_179);
  xor g141 (Z[22], n_180, n_184);
  xor g143 (n_184, A[22], B[16]);
  or g144 (n_81, wc, n_75);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_75);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_75, n_83);
endmodule

module add_signed_6_GENERIC(A, B, Z);
  input [22:0] A;
  input [16:0] B;
  output [22:0] Z;
  wire [22:0] A;
  wire [16:0] B;
  wire [22:0] Z;
  add_signed_6_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_756_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [16:0] A;
  input [18:0] B;
  output [19:0] Z;
  wire [16:0] A;
  wire [18:0] B;
  wire [19:0] Z;
  wire n_60, n_61, n_62, n_63, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154;
  not g3 (Z[19], n_61);
  nand g4 (n_63, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_68, A[1], B[1]);
  nand g13 (n_72, n_68, n_69, n_70);
  xor g14 (n_71, A[1], B[1]);
  nand g16 (n_73, A[2], B[2]);
  nand g17 (n_74, A[2], n_72);
  nand g18 (n_75, B[2], n_72);
  nand g19 (n_77, n_73, n_74, n_75);
  xor g20 (n_76, A[2], B[2]);
  xor g21 (Z[2], n_72, n_76);
  nand g22 (n_78, A[3], B[3]);
  nand g23 (n_79, A[3], n_77);
  nand g24 (n_80, B[3], n_77);
  nand g25 (n_82, n_78, n_79, n_80);
  xor g26 (n_81, A[3], B[3]);
  xor g27 (Z[3], n_77, n_81);
  nand g28 (n_83, A[4], B[4]);
  nand g29 (n_84, A[4], n_82);
  nand g30 (n_85, B[4], n_82);
  nand g31 (n_87, n_83, n_84, n_85);
  xor g32 (n_86, A[4], B[4]);
  xor g33 (Z[4], n_82, n_86);
  nand g34 (n_88, A[5], B[5]);
  nand g35 (n_89, A[5], n_87);
  nand g36 (n_90, B[5], n_87);
  nand g37 (n_92, n_88, n_89, n_90);
  xor g38 (n_91, A[5], B[5]);
  xor g39 (Z[5], n_87, n_91);
  nand g40 (n_93, A[6], B[6]);
  nand g41 (n_94, A[6], n_92);
  nand g42 (n_95, B[6], n_92);
  nand g43 (n_97, n_93, n_94, n_95);
  xor g44 (n_96, A[6], B[6]);
  xor g45 (Z[6], n_92, n_96);
  nand g46 (n_98, A[7], B[7]);
  nand g47 (n_99, A[7], n_97);
  nand g48 (n_100, B[7], n_97);
  nand g49 (n_102, n_98, n_99, n_100);
  xor g50 (n_101, A[7], B[7]);
  xor g51 (Z[7], n_97, n_101);
  nand g52 (n_60, A[8], B[8]);
  nand g53 (n_103, A[8], n_102);
  nand g54 (n_62, B[8], n_102);
  nand g55 (n_105, n_60, n_103, n_62);
  xor g56 (n_104, A[8], B[8]);
  xor g57 (Z[8], n_102, n_104);
  nand g58 (n_106, A[9], B[9]);
  nand g59 (n_107, A[9], n_105);
  nand g60 (n_108, B[9], n_105);
  nand g61 (n_110, n_106, n_107, n_108);
  xor g62 (n_109, A[9], B[9]);
  xor g63 (Z[9], n_105, n_109);
  nand g64 (n_111, A[10], B[10]);
  nand g65 (n_112, A[10], n_110);
  nand g66 (n_113, B[10], n_110);
  nand g67 (n_115, n_111, n_112, n_113);
  xor g68 (n_114, A[10], B[10]);
  xor g69 (Z[10], n_110, n_114);
  nand g70 (n_116, A[11], B[11]);
  nand g71 (n_117, A[11], n_115);
  nand g72 (n_118, B[11], n_115);
  nand g73 (n_120, n_116, n_117, n_118);
  xor g74 (n_119, A[11], B[11]);
  xor g75 (Z[11], n_115, n_119);
  nand g76 (n_121, A[12], B[12]);
  nand g77 (n_122, A[12], n_120);
  nand g78 (n_123, B[12], n_120);
  nand g79 (n_125, n_121, n_122, n_123);
  xor g80 (n_124, A[12], B[12]);
  xor g81 (Z[12], n_120, n_124);
  nand g82 (n_126, A[13], B[13]);
  nand g83 (n_127, A[13], n_125);
  nand g84 (n_128, B[13], n_125);
  nand g85 (n_130, n_126, n_127, n_128);
  xor g86 (n_129, A[13], B[13]);
  xor g87 (Z[13], n_125, n_129);
  nand g88 (n_131, A[14], B[14]);
  nand g89 (n_132, A[14], n_130);
  nand g90 (n_133, B[14], n_130);
  nand g91 (n_135, n_131, n_132, n_133);
  xor g92 (n_134, A[14], B[14]);
  xor g93 (Z[14], n_130, n_134);
  nand g94 (n_136, A[15], B[15]);
  nand g95 (n_137, A[15], n_135);
  nand g96 (n_138, B[15], n_135);
  nand g97 (n_140, n_136, n_137, n_138);
  xor g98 (n_139, A[15], B[15]);
  xor g99 (Z[15], n_135, n_139);
  nand g100 (n_141, A[16], B[16]);
  nand g101 (n_142, A[16], n_140);
  nand g102 (n_143, B[16], n_140);
  nand g103 (n_145, n_141, n_142, n_143);
  xor g104 (n_144, A[16], B[16]);
  xor g105 (Z[16], n_140, n_144);
  nand g106 (n_146, A[16], B[17]);
  nand g107 (n_147, A[16], n_145);
  nand g108 (n_148, B[17], n_145);
  nand g109 (n_150, n_146, n_147, n_148);
  xor g110 (n_149, A[16], B[17]);
  xor g111 (Z[17], n_145, n_149);
  nand g115 (n_61, n_151, n_152, n_153);
  xor g117 (Z[18], n_150, n_154);
  or g119 (n_151, A[16], B[18]);
  xor g120 (n_154, A[16], B[18]);
  or g121 (n_69, wc, n_63);
  not gc (wc, A[1]);
  or g122 (n_70, wc0, n_63);
  not gc0 (wc0, B[1]);
  xnor g123 (Z[1], n_63, n_71);
  or g124 (n_152, A[16], wc1);
  not gc1 (wc1, n_150);
  or g125 (n_153, B[18], wc2);
  not gc2 (wc2, n_150);
endmodule

module add_signed_756_GENERIC(A, B, Z);
  input [16:0] A;
  input [18:0] B;
  output [19:0] Z;
  wire [16:0] A;
  wire [18:0] B;
  wire [19:0] Z;
  add_signed_756_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_898_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [11:0] A;
  input [13:0] B;
  output [14:0] Z;
  wire [11:0] A;
  wire [13:0] B;
  wire [14:0] Z;
  wire n_45, n_46, n_47, n_48, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114;
  not g3 (Z[14], n_46);
  nand g4 (n_48, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_53, A[1], B[1]);
  nand g13 (n_57, n_53, n_54, n_55);
  xor g14 (n_56, A[1], B[1]);
  nand g16 (n_58, A[2], B[2]);
  nand g17 (n_59, A[2], n_57);
  nand g18 (n_60, B[2], n_57);
  nand g19 (n_62, n_58, n_59, n_60);
  xor g20 (n_61, A[2], B[2]);
  xor g21 (Z[2], n_57, n_61);
  nand g22 (n_63, A[3], B[3]);
  nand g23 (n_64, A[3], n_62);
  nand g24 (n_65, B[3], n_62);
  nand g25 (n_67, n_63, n_64, n_65);
  xor g26 (n_66, A[3], B[3]);
  xor g27 (Z[3], n_62, n_66);
  nand g28 (n_68, A[4], B[4]);
  nand g29 (n_69, A[4], n_67);
  nand g30 (n_70, B[4], n_67);
  nand g31 (n_72, n_68, n_69, n_70);
  xor g32 (n_71, A[4], B[4]);
  xor g33 (Z[4], n_67, n_71);
  nand g34 (n_73, A[5], B[5]);
  nand g35 (n_74, A[5], n_72);
  nand g36 (n_75, B[5], n_72);
  nand g37 (n_45, n_73, n_74, n_75);
  xor g38 (n_76, A[5], B[5]);
  xor g39 (Z[5], n_72, n_76);
  nand g40 (n_77, A[6], B[6]);
  nand g41 (n_47, A[6], n_45);
  nand g42 (n_78, B[6], n_45);
  nand g43 (n_80, n_77, n_47, n_78);
  xor g44 (n_79, A[6], B[6]);
  xor g45 (Z[6], n_45, n_79);
  nand g46 (n_81, A[7], B[7]);
  nand g47 (n_82, A[7], n_80);
  nand g48 (n_83, B[7], n_80);
  nand g49 (n_85, n_81, n_82, n_83);
  xor g50 (n_84, A[7], B[7]);
  xor g51 (Z[7], n_80, n_84);
  nand g52 (n_86, A[8], B[8]);
  nand g53 (n_87, A[8], n_85);
  nand g54 (n_88, B[8], n_85);
  nand g55 (n_90, n_86, n_87, n_88);
  xor g56 (n_89, A[8], B[8]);
  xor g57 (Z[8], n_85, n_89);
  nand g58 (n_91, A[9], B[9]);
  nand g59 (n_92, A[9], n_90);
  nand g60 (n_93, B[9], n_90);
  nand g61 (n_95, n_91, n_92, n_93);
  xor g62 (n_94, A[9], B[9]);
  xor g63 (Z[9], n_90, n_94);
  nand g64 (n_96, A[10], B[10]);
  nand g65 (n_97, A[10], n_95);
  nand g66 (n_98, B[10], n_95);
  nand g67 (n_100, n_96, n_97, n_98);
  xor g68 (n_99, A[10], B[10]);
  xor g69 (Z[10], n_95, n_99);
  nand g70 (n_101, A[11], B[11]);
  nand g71 (n_102, A[11], n_100);
  nand g72 (n_103, B[11], n_100);
  nand g73 (n_105, n_101, n_102, n_103);
  xor g74 (n_104, A[11], B[11]);
  xor g75 (Z[11], n_100, n_104);
  nand g76 (n_106, A[11], B[12]);
  nand g77 (n_107, A[11], n_105);
  nand g78 (n_108, B[12], n_105);
  nand g79 (n_110, n_106, n_107, n_108);
  xor g80 (n_109, A[11], B[12]);
  xor g81 (Z[12], n_105, n_109);
  nand g85 (n_46, n_111, n_112, n_113);
  xor g87 (Z[13], n_110, n_114);
  or g89 (n_111, A[11], B[13]);
  xor g90 (n_114, A[11], B[13]);
  or g91 (n_54, wc, n_48);
  not gc (wc, A[1]);
  or g92 (n_55, wc0, n_48);
  not gc0 (wc0, B[1]);
  xnor g93 (Z[1], n_48, n_56);
  or g94 (n_112, A[11], wc1);
  not gc1 (wc1, n_110);
  or g95 (n_113, B[13], wc2);
  not gc2 (wc2, n_110);
endmodule

module add_signed_898_GENERIC(A, B, Z);
  input [11:0] A;
  input [13:0] B;
  output [14:0] Z;
  wire [11:0] A;
  wire [13:0] B;
  wire [14:0] Z;
  add_signed_898_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module increment_unsigned_752_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [17:0] A;
  input CI;
  output [17:0] Z;
  wire [17:0] A;
  wire CI;
  wire [17:0] Z;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_38, A[0], CI);
  xor g18 (Z[1], A[1], n_38);
  and g19 (n_39, A[1], n_38);
  xor g20 (Z[2], A[2], n_39);
  and g21 (n_40, A[2], n_39);
  xor g22 (Z[3], A[3], n_40);
  and g23 (n_41, A[3], n_40);
  xor g24 (Z[4], A[4], n_41);
  and g25 (n_42, A[4], n_41);
  xor g26 (Z[5], A[5], n_42);
  and g27 (n_43, A[5], n_42);
  xor g28 (Z[6], A[6], n_43);
  and g29 (n_44, A[6], n_43);
  xor g30 (Z[7], A[7], n_44);
  and g31 (n_45, A[7], n_44);
  xor g32 (Z[8], A[8], n_45);
  and g33 (n_46, A[8], n_45);
  xor g34 (Z[9], A[9], n_46);
  and g35 (n_47, A[9], n_46);
  xor g36 (Z[10], A[10], n_47);
  and g37 (n_48, A[10], n_47);
  xor g38 (Z[11], A[11], n_48);
  and g39 (n_49, A[11], n_48);
  xor g40 (Z[12], A[12], n_49);
  and g41 (n_50, A[12], n_49);
  xor g42 (Z[13], A[13], n_50);
  and g43 (n_51, A[13], n_50);
  xor g44 (Z[14], A[14], n_51);
  and g45 (n_52, A[14], n_51);
  xor g46 (Z[15], A[15], n_52);
  and g47 (n_53, A[15], n_52);
  xor g48 (Z[16], A[16], n_53);
  and g49 (n_54, A[16], n_53);
  xor g50 (Z[17], A[17], n_54);
endmodule

module increment_unsigned_752_GENERIC(A, CI, Z);
  input [17:0] A;
  input CI;
  output [17:0] Z;
  wire [17:0] A;
  wire CI;
  wire [17:0] Z;
  increment_unsigned_752_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_752_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [17:0] A;
  input CI;
  output [17:0] Z;
  wire [17:0] A;
  wire CI;
  wire [17:0] Z;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_38, A[0], CI);
  xor g18 (Z[1], A[1], n_38);
  and g19 (n_39, A[1], n_38);
  xor g20 (Z[2], A[2], n_39);
  and g21 (n_40, A[2], n_39);
  xor g22 (Z[3], A[3], n_40);
  and g23 (n_41, A[3], n_40);
  xor g24 (Z[4], A[4], n_41);
  and g25 (n_42, A[4], n_41);
  xor g26 (Z[5], A[5], n_42);
  and g27 (n_43, A[5], n_42);
  xor g28 (Z[6], A[6], n_43);
  and g29 (n_44, A[6], n_43);
  xor g30 (Z[7], A[7], n_44);
  and g31 (n_45, A[7], n_44);
  xor g32 (Z[8], A[8], n_45);
  and g33 (n_46, A[8], n_45);
  xor g34 (Z[9], A[9], n_46);
  and g35 (n_47, A[9], n_46);
  xor g36 (Z[10], A[10], n_47);
  and g37 (n_48, A[10], n_47);
  xor g38 (Z[11], A[11], n_48);
  and g39 (n_49, A[11], n_48);
  xor g40 (Z[12], A[12], n_49);
  and g41 (n_50, A[12], n_49);
  xor g42 (Z[13], A[13], n_50);
  and g43 (n_51, A[13], n_50);
  xor g44 (Z[14], A[14], n_51);
  and g45 (n_52, A[14], n_51);
  xor g46 (Z[15], A[15], n_52);
  and g47 (n_53, A[15], n_52);
  xor g48 (Z[16], A[16], n_53);
  and g49 (n_54, A[16], n_53);
  xor g50 (Z[17], A[17], n_54);
endmodule

module increment_unsigned_752_1_GENERIC(A, CI, Z);
  input [17:0] A;
  input CI;
  output [17:0] Z;
  wire [17:0] A;
  wire CI;
  wire [17:0] Z;
  increment_unsigned_752_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_753_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [21:0] A;
  input CI;
  output [21:0] Z;
  wire [21:0] A;
  wire CI;
  wire [21:0] Z;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_46, A[0], CI);
  xor g22 (Z[1], A[1], n_46);
  and g23 (n_47, A[1], n_46);
  xor g24 (Z[2], A[2], n_47);
  and g25 (n_48, A[2], n_47);
  xor g26 (Z[3], A[3], n_48);
  and g27 (n_49, A[3], n_48);
  xor g28 (Z[4], A[4], n_49);
  and g29 (n_50, A[4], n_49);
  xor g30 (Z[5], A[5], n_50);
  and g31 (n_51, A[5], n_50);
  xor g32 (Z[6], A[6], n_51);
  and g33 (n_52, A[6], n_51);
  xor g34 (Z[7], A[7], n_52);
  and g35 (n_53, A[7], n_52);
  xor g36 (Z[8], A[8], n_53);
  and g37 (n_54, A[8], n_53);
  xor g38 (Z[9], A[9], n_54);
  and g39 (n_55, A[9], n_54);
  xor g40 (Z[10], A[10], n_55);
  and g41 (n_56, A[10], n_55);
  xor g42 (Z[11], A[11], n_56);
  and g43 (n_57, A[11], n_56);
  xor g44 (Z[12], A[12], n_57);
  and g45 (n_58, A[12], n_57);
  xor g46 (Z[13], A[13], n_58);
  and g47 (n_59, A[13], n_58);
  xor g48 (Z[14], A[14], n_59);
  and g49 (n_60, A[14], n_59);
  xor g50 (Z[15], A[15], n_60);
  and g51 (n_61, A[15], n_60);
  xor g52 (Z[16], A[16], n_61);
  and g53 (n_62, A[16], n_61);
  xor g54 (Z[17], A[17], n_62);
  and g55 (n_63, A[17], n_62);
  xor g56 (Z[18], A[18], n_63);
  and g57 (n_64, A[18], n_63);
  xor g58 (Z[19], A[19], n_64);
  and g59 (n_65, A[19], n_64);
  xor g60 (Z[20], A[20], n_65);
  and g61 (n_66, A[20], n_65);
  xor g62 (Z[21], A[21], n_66);
endmodule

module increment_unsigned_753_GENERIC(A, CI, Z);
  input [21:0] A;
  input CI;
  output [21:0] Z;
  wire [21:0] A;
  wire CI;
  wire [21:0] Z;
  increment_unsigned_753_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_753_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [21:0] A;
  input CI;
  output [21:0] Z;
  wire [21:0] A;
  wire CI;
  wire [21:0] Z;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_46, A[0], CI);
  xor g22 (Z[1], A[1], n_46);
  and g23 (n_47, A[1], n_46);
  xor g24 (Z[2], A[2], n_47);
  and g25 (n_48, A[2], n_47);
  xor g26 (Z[3], A[3], n_48);
  and g27 (n_49, A[3], n_48);
  xor g28 (Z[4], A[4], n_49);
  and g29 (n_50, A[4], n_49);
  xor g30 (Z[5], A[5], n_50);
  and g31 (n_51, A[5], n_50);
  xor g32 (Z[6], A[6], n_51);
  and g33 (n_52, A[6], n_51);
  xor g34 (Z[7], A[7], n_52);
  and g35 (n_53, A[7], n_52);
  xor g36 (Z[8], A[8], n_53);
  and g37 (n_54, A[8], n_53);
  xor g38 (Z[9], A[9], n_54);
  and g39 (n_55, A[9], n_54);
  xor g40 (Z[10], A[10], n_55);
  and g41 (n_56, A[10], n_55);
  xor g42 (Z[11], A[11], n_56);
  and g43 (n_57, A[11], n_56);
  xor g44 (Z[12], A[12], n_57);
  and g45 (n_58, A[12], n_57);
  xor g46 (Z[13], A[13], n_58);
  and g47 (n_59, A[13], n_58);
  xor g48 (Z[14], A[14], n_59);
  and g49 (n_60, A[14], n_59);
  xor g50 (Z[15], A[15], n_60);
  and g51 (n_61, A[15], n_60);
  xor g52 (Z[16], A[16], n_61);
  and g53 (n_62, A[16], n_61);
  xor g54 (Z[17], A[17], n_62);
  and g55 (n_63, A[17], n_62);
  xor g56 (Z[18], A[18], n_63);
  and g57 (n_64, A[18], n_63);
  xor g58 (Z[19], A[19], n_64);
  and g59 (n_65, A[19], n_64);
  xor g60 (Z[20], A[20], n_65);
  and g61 (n_66, A[20], n_65);
  xor g62 (Z[21], A[21], n_66);
endmodule

module increment_unsigned_753_1_GENERIC(A, CI, Z);
  input [21:0] A;
  input CI;
  output [21:0] Z;
  wire [21:0] A;
  wire CI;
  wire [21:0] Z;
  increment_unsigned_753_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_755_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_36, A[0], CI);
  xor g17 (Z[1], A[1], n_36);
  and g18 (n_37, A[1], n_36);
  xor g19 (Z[2], A[2], n_37);
  and g20 (n_38, A[2], n_37);
  xor g21 (Z[3], A[3], n_38);
  and g22 (n_39, A[3], n_38);
  xor g23 (Z[4], A[4], n_39);
  and g24 (n_40, A[4], n_39);
  xor g25 (Z[5], A[5], n_40);
  and g26 (n_41, A[5], n_40);
  xor g27 (Z[6], A[6], n_41);
  and g28 (n_42, A[6], n_41);
  xor g29 (Z[7], A[7], n_42);
  and g30 (n_43, A[7], n_42);
  xor g31 (Z[8], A[8], n_43);
  and g32 (n_44, A[8], n_43);
  xor g33 (Z[9], A[9], n_44);
  and g34 (n_45, A[9], n_44);
  xor g35 (Z[10], A[10], n_45);
  and g36 (n_46, A[10], n_45);
  xor g37 (Z[11], A[11], n_46);
  and g38 (n_47, A[11], n_46);
  xor g39 (Z[12], A[12], n_47);
  and g40 (n_48, A[12], n_47);
  xor g41 (Z[13], A[13], n_48);
  and g42 (n_49, A[13], n_48);
  xor g43 (Z[14], A[14], n_49);
  and g44 (n_50, A[14], n_49);
  xor g45 (Z[15], A[15], n_50);
  and g46 (n_51, A[15], n_50);
  xor g47 (Z[16], A[16], n_51);
endmodule

module increment_unsigned_755_GENERIC(A, CI, Z);
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  increment_unsigned_755_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_755_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_36, A[0], CI);
  xor g17 (Z[1], A[1], n_36);
  and g18 (n_37, A[1], n_36);
  xor g19 (Z[2], A[2], n_37);
  and g20 (n_38, A[2], n_37);
  xor g21 (Z[3], A[3], n_38);
  and g22 (n_39, A[3], n_38);
  xor g23 (Z[4], A[4], n_39);
  and g24 (n_40, A[4], n_39);
  xor g25 (Z[5], A[5], n_40);
  and g26 (n_41, A[5], n_40);
  xor g27 (Z[6], A[6], n_41);
  and g28 (n_42, A[6], n_41);
  xor g29 (Z[7], A[7], n_42);
  and g30 (n_43, A[7], n_42);
  xor g31 (Z[8], A[8], n_43);
  and g32 (n_44, A[8], n_43);
  xor g33 (Z[9], A[9], n_44);
  and g34 (n_45, A[9], n_44);
  xor g35 (Z[10], A[10], n_45);
  and g36 (n_46, A[10], n_45);
  xor g37 (Z[11], A[11], n_46);
  and g38 (n_47, A[11], n_46);
  xor g39 (Z[12], A[12], n_47);
  and g40 (n_48, A[12], n_47);
  xor g41 (Z[13], A[13], n_48);
  and g42 (n_49, A[13], n_48);
  xor g43 (Z[14], A[14], n_49);
  and g44 (n_50, A[14], n_49);
  xor g45 (Z[15], A[15], n_50);
  and g46 (n_51, A[15], n_50);
  xor g47 (Z[16], A[16], n_51);
endmodule

module increment_unsigned_755_1_GENERIC(A, CI, Z);
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  increment_unsigned_755_1_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_755_2_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_36, A[0], CI);
  xor g17 (Z[1], A[1], n_36);
  and g18 (n_37, A[1], n_36);
  xor g19 (Z[2], A[2], n_37);
  and g20 (n_38, A[2], n_37);
  xor g21 (Z[3], A[3], n_38);
  and g22 (n_39, A[3], n_38);
  xor g23 (Z[4], A[4], n_39);
  and g24 (n_40, A[4], n_39);
  xor g25 (Z[5], A[5], n_40);
  and g26 (n_41, A[5], n_40);
  xor g27 (Z[6], A[6], n_41);
  and g28 (n_42, A[6], n_41);
  xor g29 (Z[7], A[7], n_42);
  and g30 (n_43, A[7], n_42);
  xor g31 (Z[8], A[8], n_43);
  and g32 (n_44, A[8], n_43);
  xor g33 (Z[9], A[9], n_44);
  and g34 (n_45, A[9], n_44);
  xor g35 (Z[10], A[10], n_45);
  and g36 (n_46, A[10], n_45);
  xor g37 (Z[11], A[11], n_46);
  and g38 (n_47, A[11], n_46);
  xor g39 (Z[12], A[12], n_47);
  and g40 (n_48, A[12], n_47);
  xor g41 (Z[13], A[13], n_48);
  and g42 (n_49, A[13], n_48);
  xor g43 (Z[14], A[14], n_49);
  and g44 (n_50, A[14], n_49);
  xor g45 (Z[15], A[15], n_50);
  and g46 (n_51, A[15], n_50);
  xor g47 (Z[16], A[16], n_51);
endmodule

module increment_unsigned_755_2_GENERIC(A, CI, Z);
  input [16:0] A;
  input CI;
  output [16:0] Z;
  wire [16:0] A;
  wire CI;
  wire [16:0] Z;
  increment_unsigned_755_2_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_762_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_40, A[0], CI);
  xor g19 (Z[1], A[1], n_40);
  and g20 (n_41, A[1], n_40);
  xor g21 (Z[2], A[2], n_41);
  and g22 (n_42, A[2], n_41);
  xor g23 (Z[3], A[3], n_42);
  and g24 (n_43, A[3], n_42);
  xor g25 (Z[4], A[4], n_43);
  and g26 (n_44, A[4], n_43);
  xor g27 (Z[5], A[5], n_44);
  and g28 (n_45, A[5], n_44);
  xor g29 (Z[6], A[6], n_45);
  and g30 (n_46, A[6], n_45);
  xor g31 (Z[7], A[7], n_46);
  and g32 (n_47, A[7], n_46);
  xor g33 (Z[8], A[8], n_47);
  and g34 (n_48, A[8], n_47);
  xor g35 (Z[9], A[9], n_48);
  and g36 (n_49, A[9], n_48);
  xor g37 (Z[10], A[10], n_49);
  and g38 (n_50, A[10], n_49);
  xor g39 (Z[11], A[11], n_50);
  and g40 (n_51, A[11], n_50);
  xor g41 (Z[12], A[12], n_51);
  and g42 (n_52, A[12], n_51);
  xor g43 (Z[13], A[13], n_52);
  and g44 (n_53, A[13], n_52);
  xor g45 (Z[14], A[14], n_53);
  and g46 (n_54, A[14], n_53);
  xor g47 (Z[15], A[15], n_54);
  and g48 (n_55, A[15], n_54);
  xor g49 (Z[16], A[16], n_55);
  and g50 (n_56, A[16], n_55);
  xor g51 (Z[17], A[17], n_56);
  and g52 (n_57, A[17], n_56);
  xor g53 (Z[18], A[18], n_57);
endmodule

module increment_unsigned_762_GENERIC(A, CI, Z);
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  increment_unsigned_762_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module mult_signed_const_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * -209;"
  input [16:0] A;
  output [25:0] Z;
  wire [16:0] A;
  wire [25:0] Z;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_43, n_46, n_47, n_48, n_49, n_50, n_51;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_102, n_105, n_106;
  wire n_107, n_109, n_110, n_111, n_112, n_114, n_115, n_116;
  wire n_117, n_119, n_120, n_121, n_123, n_124, n_125, n_126;
  wire n_128, n_129, n_130, n_131, n_133, n_134, n_135, n_136;
  wire n_138, n_139, n_140, n_141, n_143, n_144, n_145, n_146;
  wire n_148, n_149, n_150, n_151, n_153, n_154, n_155, n_156;
  wire n_158, n_159, n_160, n_161, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_171, n_172, n_173, n_176, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_256, n_258, n_259, n_260, n_261, n_264, n_266, n_267;
  wire n_268, n_269, n_272, n_274, n_275, n_276, n_277, n_280;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_296, n_298, n_299, n_300;
  wire n_301, n_315, n_320, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  assign Z[0] = A[0];
  assign Z[24] = Z[25];
  xor g72 (n_63, A[0], n_102);
  nand g84 (n_111, A[0], A[1], n_181);
  xor g85 (n_182, n_105, n_106);
  xor g86 (n_62, n_182, n_107);
  nand g87 (n_183, n_105, n_106);
  nand g88 (n_184, n_107, n_106);
  nand g89 (n_185, n_105, n_107);
  nand g90 (n_35, n_183, n_184, n_185);
  xor g94 (n_112, n_186, n_109);
  nand g98 (n_117, n_187, n_188, n_189);
  xor g99 (n_190, n_110, n_111);
  xor g100 (n_61, n_190, n_112);
  nand g101 (n_191, n_110, n_111);
  nand g102 (n_192, n_112, n_111);
  nand g103 (n_193, n_110, n_112);
  nand g104 (n_34, n_191, n_192, n_193);
  xor g108 (n_116, n_194, n_114);
  nand g112 (n_121, n_195, n_196, n_197);
  xor g113 (n_198, n_115, n_116);
  xor g114 (n_60, n_198, n_117);
  nand g115 (n_199, n_115, n_116);
  nand g116 (n_200, n_117, n_116);
  nand g117 (n_201, n_115, n_117);
  nand g118 (n_33, n_199, n_200, n_201);
  xor g122 (n_120, n_202, n_43);
  nand g126 (n_126, n_203, n_204, n_205);
  xor g127 (n_206, n_119, n_120);
  xor g128 (n_59, n_206, n_121);
  nand g129 (n_207, n_119, n_120);
  nand g130 (n_208, n_121, n_120);
  nand g131 (n_209, n_119, n_121);
  nand g132 (n_32, n_207, n_208, n_209);
  xor g136 (n_125, n_210, n_123);
  nand g140 (n_131, n_211, n_212, n_213);
  xor g141 (n_214, n_124, n_125);
  xor g142 (n_58, n_214, n_126);
  nand g143 (n_215, n_124, n_125);
  nand g144 (n_216, n_126, n_125);
  nand g145 (n_217, n_124, n_126);
  nand g146 (n_31, n_215, n_216, n_217);
  xor g150 (n_130, n_218, n_128);
  nand g154 (n_136, n_219, n_220, n_221);
  xor g155 (n_222, n_129, n_130);
  xor g156 (n_57, n_222, n_131);
  nand g157 (n_223, n_129, n_130);
  nand g158 (n_224, n_131, n_130);
  nand g159 (n_225, n_129, n_131);
  nand g160 (n_30, n_223, n_224, n_225);
  xor g164 (n_135, n_226, n_133);
  nand g168 (n_141, n_227, n_228, n_229);
  xor g169 (n_230, n_134, n_135);
  xor g170 (n_56, n_230, n_136);
  nand g171 (n_231, n_134, n_135);
  nand g172 (n_232, n_136, n_135);
  nand g173 (n_233, n_134, n_136);
  nand g174 (n_29, n_231, n_232, n_233);
  xor g178 (n_140, n_234, n_138);
  nand g182 (n_146, n_235, n_236, n_237);
  xor g183 (n_238, n_139, n_140);
  xor g184 (n_55, n_238, n_141);
  nand g185 (n_239, n_139, n_140);
  nand g186 (n_240, n_141, n_140);
  nand g187 (n_241, n_139, n_141);
  nand g188 (n_28, n_239, n_240, n_241);
  xor g192 (n_145, n_242, n_143);
  nand g196 (n_151, n_243, n_244, n_245);
  xor g197 (n_246, n_144, n_145);
  xor g198 (n_54, n_246, n_146);
  nand g199 (n_247, n_144, n_145);
  nand g200 (n_248, n_146, n_145);
  nand g201 (n_249, n_144, n_146);
  nand g202 (n_27, n_247, n_248, n_249);
  nand g208 (n_154, n_251, n_252, n_253);
  xor g210 (n_150, A[10], n_148);
  xor g215 (n_258, n_149, n_150);
  xor g216 (n_53, n_258, n_151);
  nand g217 (n_259, n_149, n_150);
  nand g218 (n_260, n_151, n_150);
  nand g219 (n_261, n_149, n_151);
  nand g220 (n_26, n_259, n_260, n_261);
  xor g224 (n_155, A[10], n_153);
  xor g229 (n_266, n_154, n_155);
  xor g230 (n_52, n_266, n_156);
  nand g231 (n_267, n_154, n_155);
  nand g232 (n_268, n_156, n_155);
  nand g233 (n_269, n_154, n_156);
  nand g234 (n_25, n_267, n_268, n_269);
  xor g238 (n_160, A[11], n_158);
  xor g243 (n_274, n_159, n_160);
  xor g244 (n_51, n_274, n_161);
  nand g245 (n_275, n_159, n_160);
  nand g246 (n_276, n_161, n_160);
  nand g247 (n_277, n_159, n_161);
  nand g248 (n_24, n_275, n_276, n_277);
  xor g252 (n_165, A[12], n_163);
  xor g257 (n_282, n_164, n_165);
  xor g258 (n_50, n_282, n_166);
  nand g259 (n_283, n_164, n_165);
  nand g260 (n_284, n_166, n_165);
  nand g261 (n_285, n_164, n_166);
  nand g262 (n_23, n_283, n_284, n_285);
  nand g268 (n_172, n_287, n_288, n_289);
  xor g269 (n_290, n_167, n_168);
  xor g270 (n_49, n_290, n_169);
  nand g271 (n_291, n_167, n_168);
  nand g272 (n_292, n_169, n_168);
  nand g273 (n_293, n_167, n_169);
  nand g274 (n_48, n_291, n_292, n_293);
  nand g280 (n_296, n_172, n_171);
  xor g284 (n_21, n_298, n_173);
  nand g287 (n_301, A[16], n_173);
  nand g288 (n_46, n_299, n_300, n_301);
  nand g31 (n_328, n_324, n_325, n_326);
  nand g36 (n_331, n_64, n_328);
  nand g37 (n_333, n_329, n_330, n_331);
  xor g39 (Z[5], n_328, n_332);
  nand g40 (n_334, n_37, n_63);
  nand g41 (n_335, n_37, n_333);
  nand g42 (n_336, n_63, n_333);
  nand g43 (n_338, n_334, n_335, n_336);
  xor g44 (n_337, n_37, n_63);
  xor g45 (Z[6], n_333, n_337);
  nand g46 (n_339, n_36, n_62);
  nand g47 (n_340, n_36, n_338);
  nand g48 (n_341, n_62, n_338);
  nand g49 (n_343, n_339, n_340, n_341);
  xor g50 (n_342, n_36, n_62);
  xor g51 (Z[7], n_338, n_342);
  nand g52 (n_344, n_35, n_61);
  nand g53 (n_345, n_35, n_343);
  nand g54 (n_346, n_61, n_343);
  nand g55 (n_348, n_344, n_345, n_346);
  xor g56 (n_347, n_35, n_61);
  xor g57 (Z[8], n_343, n_347);
  nand g58 (n_349, n_34, n_60);
  nand g59 (n_350, n_34, n_348);
  nand g60 (n_351, n_60, n_348);
  nand g61 (n_353, n_349, n_350, n_351);
  xor g62 (n_352, n_34, n_60);
  xor g63 (Z[9], n_348, n_352);
  nand g64 (n_354, n_33, n_59);
  nand g304 (n_355, n_33, n_353);
  nand g305 (n_356, n_59, n_353);
  nand g306 (n_358, n_354, n_355, n_356);
  xor g307 (n_357, n_33, n_59);
  xor g308 (Z[10], n_353, n_357);
  nand g309 (n_359, n_32, n_58);
  nand g310 (n_360, n_32, n_358);
  nand g311 (n_361, n_58, n_358);
  nand g312 (n_363, n_359, n_360, n_361);
  xor g313 (n_362, n_32, n_58);
  xor g314 (Z[11], n_358, n_362);
  nand g315 (n_364, n_31, n_57);
  nand g316 (n_365, n_31, n_363);
  nand g317 (n_366, n_57, n_363);
  nand g318 (n_368, n_364, n_365, n_366);
  xor g319 (n_367, n_31, n_57);
  xor g320 (Z[12], n_363, n_367);
  nand g321 (n_369, n_30, n_56);
  nand g322 (n_370, n_30, n_368);
  nand g323 (n_371, n_56, n_368);
  nand g324 (n_373, n_369, n_370, n_371);
  xor g325 (n_372, n_30, n_56);
  xor g326 (Z[13], n_368, n_372);
  nand g327 (n_374, n_29, n_55);
  nand g328 (n_375, n_29, n_373);
  nand g329 (n_376, n_55, n_373);
  nand g330 (n_378, n_374, n_375, n_376);
  xor g331 (n_377, n_29, n_55);
  xor g332 (Z[14], n_373, n_377);
  nand g333 (n_379, n_28, n_54);
  nand g334 (n_380, n_28, n_378);
  nand g335 (n_381, n_54, n_378);
  nand g336 (n_383, n_379, n_380, n_381);
  xor g337 (n_382, n_28, n_54);
  xor g338 (Z[15], n_378, n_382);
  nand g339 (n_384, n_27, n_53);
  nand g340 (n_385, n_27, n_383);
  nand g341 (n_386, n_53, n_383);
  nand g342 (n_388, n_384, n_385, n_386);
  xor g343 (n_387, n_27, n_53);
  xor g344 (Z[16], n_383, n_387);
  nand g345 (n_389, n_26, n_52);
  nand g346 (n_390, n_26, n_388);
  nand g347 (n_391, n_52, n_388);
  nand g348 (n_393, n_389, n_390, n_391);
  xor g349 (n_392, n_26, n_52);
  xor g350 (Z[17], n_388, n_392);
  nand g351 (n_394, n_25, n_51);
  nand g352 (n_395, n_25, n_393);
  nand g353 (n_396, n_51, n_393);
  nand g354 (n_398, n_394, n_395, n_396);
  xor g355 (n_397, n_25, n_51);
  xor g356 (Z[18], n_393, n_397);
  nand g357 (n_399, n_24, n_50);
  nand g358 (n_400, n_24, n_398);
  nand g359 (n_401, n_50, n_398);
  nand g360 (n_403, n_399, n_400, n_401);
  xor g361 (n_402, n_24, n_50);
  xor g362 (Z[19], n_398, n_402);
  nand g363 (n_404, n_23, n_49);
  nand g364 (n_405, n_23, n_403);
  nand g365 (n_406, n_49, n_403);
  nand g366 (n_408, n_404, n_405, n_406);
  xor g367 (n_407, n_23, n_49);
  xor g368 (Z[20], n_403, n_407);
  nand g369 (n_409, n_22, n_48);
  nand g370 (n_410, n_22, n_408);
  nand g371 (n_411, n_48, n_408);
  nand g372 (n_413, n_409, n_410, n_411);
  xor g373 (n_412, n_22, n_48);
  xor g374 (Z[21], n_408, n_412);
  nand g375 (n_414, n_21, n_47);
  nand g376 (n_415, n_21, n_413);
  nand g377 (n_416, n_47, n_413);
  nand g378 (n_418, n_414, n_415, n_416);
  xor g379 (n_417, n_21, n_47);
  xor g380 (Z[22], n_413, n_417);
  nand g381 (n_419, A[16], n_46);
  nand g382 (n_420, A[16], n_418);
  nand g383 (n_421, n_46, n_418);
  nand g384 (n_423, n_419, n_420, n_421);
  xor g385 (n_422, A[16], n_46);
  xor g386 (Z[23], n_418, n_422);
  xor g395 (n_64, A[5], A[1]);
  nor g396 (n_37, A[5], A[1]);
  xor g397 (n_102, A[6], A[2]);
  nor g398 (n_106, A[6], A[2]);
  xor g399 (n_105, A[7], A[3]);
  nor g400 (n_109, A[7], A[3]);
  or g401 (n_181, A[1], A[0]);
  xor g402 (n_110, A[8], A[4]);
  nor g403 (n_114, A[8], A[4]);
  xor g404 (n_186, A[2], A[1]);
  or g405 (n_187, A[2], A[1]);
  xor g406 (n_115, A[9], A[5]);
  nor g407 (n_43, A[9], A[5]);
  xor g408 (n_194, A[3], A[2]);
  or g409 (n_195, A[3], A[2]);
  xor g410 (n_119, A[10], A[6]);
  nor g411 (n_123, A[10], A[6]);
  xor g412 (n_202, A[4], A[3]);
  or g413 (n_203, A[4], A[3]);
  xor g414 (n_124, A[11], A[7]);
  nor g415 (n_128, A[11], A[7]);
  xor g416 (n_210, A[5], A[4]);
  or g417 (n_211, A[5], A[4]);
  xor g418 (n_129, A[12], A[8]);
  nor g419 (n_133, A[12], A[8]);
  xor g420 (n_218, A[6], A[5]);
  or g421 (n_219, A[6], A[5]);
  xor g422 (n_134, A[13], A[9]);
  nor g423 (n_138, A[13], A[9]);
  xor g424 (n_226, A[7], A[6]);
  or g425 (n_227, A[7], A[6]);
  xor g426 (n_139, A[14], A[10]);
  nor g427 (n_143, A[14], A[10]);
  xor g428 (n_234, A[8], A[7]);
  or g429 (n_235, A[8], A[7]);
  xor g430 (n_144, A[15], A[11]);
  nor g431 (n_148, A[15], A[11]);
  xor g432 (n_242, A[9], A[8]);
  or g433 (n_243, A[9], A[8]);
  xnor g434 (n_250, A[16], A[12]);
  or g435 (n_251, A[12], wc);
  not gc (wc, A[16]);
  or g436 (n_252, A[12], A[9]);
  or g437 (n_253, A[9], wc0);
  not gc0 (wc0, A[16]);
  xor g438 (n_153, A[13], A[11]);
  nor g439 (n_158, A[13], A[11]);
  xor g440 (n_159, A[14], A[12]);
  nor g441 (n_163, A[14], A[12]);
  xor g442 (n_164, A[15], A[13]);
  nor g443 (n_167, A[15], A[13]);
  xnor g444 (n_286, A[16], A[14]);
  or g445 (n_287, A[14], wc1);
  not gc1 (wc1, A[16]);
  or g446 (n_288, A[14], A[13]);
  or g447 (n_289, A[13], wc2);
  not gc2 (wc2, A[16]);
  xor g448 (n_171, A[15], A[14]);
  nor g449 (n_173, A[15], A[14]);
  xnor g450 (n_298, A[16], A[15]);
  or g451 (n_299, A[15], wc3);
  not gc3 (wc3, A[16]);
  or g452 (n_176, A[0], wc4);
  not gc4 (wc4, n_102);
  xnor g454 (n_107, A[1], A[0]);
  or g455 (n_188, A[2], wc5);
  not gc5 (wc5, n_109);
  or g456 (n_189, A[1], wc6);
  not gc6 (wc6, n_109);
  or g457 (n_196, A[3], wc7);
  not gc7 (wc7, n_114);
  or g458 (n_197, A[2], wc8);
  not gc8 (wc8, n_114);
  or g459 (n_204, A[4], wc9);
  not gc9 (wc9, n_43);
  or g460 (n_205, A[3], wc10);
  not gc10 (wc10, n_43);
  or g461 (n_212, A[5], wc11);
  not gc11 (wc11, n_123);
  or g462 (n_213, A[4], wc12);
  not gc12 (wc12, n_123);
  or g463 (n_220, A[6], wc13);
  not gc13 (wc13, n_128);
  or g464 (n_221, A[5], wc14);
  not gc14 (wc14, n_128);
  or g465 (n_228, A[7], wc15);
  not gc15 (wc15, n_133);
  or g466 (n_229, A[6], wc16);
  not gc16 (wc16, n_133);
  or g467 (n_236, A[8], wc17);
  not gc17 (wc17, n_138);
  or g468 (n_237, A[7], wc18);
  not gc18 (wc18, n_138);
  or g469 (n_244, A[9], wc19);
  not gc19 (wc19, n_143);
  or g470 (n_245, A[8], wc20);
  not gc20 (wc20, n_143);
  xnor g471 (n_149, n_250, A[9]);
  or g472 (n_256, A[10], wc21);
  not gc21 (wc21, n_148);
  or g474 (n_264, A[10], wc22);
  not gc22 (wc22, n_153);
  or g476 (n_272, A[11], wc23);
  not gc23 (wc23, n_158);
  or g478 (n_280, A[12], wc24);
  not gc24 (wc24, n_163);
  xnor g480 (n_168, n_286, A[13]);
  or g482 (n_300, A[15], wc25);
  not gc25 (wc25, n_173);
  or g483 (n_324, A[0], wc26);
  not gc26 (wc26, A[4]);
  xnor g484 (n_327, A[4], A[0]);
  or g485 (n_329, A[4], wc27);
  not gc27 (wc27, n_64);
  xnor g486 (n_332, n_64, A[4]);
  or g487 (n_36, wc28, wc29, n_102);
  not gc29 (wc29, n_176);
  not gc28 (wc28, A[0]);
  or g488 (n_156, wc30, wc31, n_148);
  not gc31 (wc31, n_256);
  not gc30 (wc30, A[10]);
  or g489 (n_161, wc32, wc33, n_153);
  not gc33 (wc33, n_264);
  not gc32 (wc32, A[10]);
  or g490 (n_166, wc34, wc35, n_158);
  not gc35 (wc35, n_272);
  not gc34 (wc34, A[11]);
  or g491 (n_169, wc36, wc37, n_163);
  not gc37 (wc37, n_280);
  not gc36 (wc36, A[12]);
  xnor g492 (n_22, n_172, n_171);
  not g494 (Z[1], n_107);
  or g495 (n_47, n_171, wc38, n_172);
  not gc38 (wc38, n_296);
  or g497 (n_315, n_181, A[2]);
  xor g498 (Z[2], n_181, A[2]);
  or g500 (n_320, n_315, A[3]);
  xor g501 (Z[3], n_315, A[3]);
  or g503 (n_325, n_320, A[0]);
  or g504 (n_326, wc39, n_320);
  not gc39 (wc39, A[4]);
  xnor g505 (Z[4], n_327, n_320);
  or g506 (n_330, A[4], wc40);
  not gc40 (wc40, n_328);
  not g507 (Z[25], n_423);
endmodule

module mult_signed_const_GENERIC(A, Z);
  input [16:0] A;
  output [25:0] Z;
  wire [16:0] A;
  wire [25:0] Z;
  mult_signed_const_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_107_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 209;"
  input [16:0] A;
  output [24:0] Z;
  wire [16:0] A;
  wire [24:0] Z;
  wire n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27;
  wire n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35;
  wire n_37, n_38, n_39, n_41, n_42, n_44, n_45, n_46;
  wire n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_114, n_115, n_116, n_117, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_201, n_202, n_203, n_204;
  wire n_205, n_208, n_210, n_211, n_212, n_213, n_216, n_218;
  wire n_219, n_220, n_221, n_224, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_240, n_242, n_243, n_244, n_245, n_268, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  assign Z[2] = A[2];
  assign Z[3] = A[3];
  xor g38 (n_61, A[6], A[0]);
  and g2 (n_35, A[6], A[0]);
  xor g39 (n_94, A[7], A[3]);
  and g40 (n_95, A[7], A[3]);
  xor g41 (n_130, A[0], A[1]);
  xor g42 (n_60, n_130, n_94);
  nand g3 (n_131, A[0], A[1]);
  nand g4 (n_132, n_94, A[1]);
  nand g43 (n_133, A[0], n_94);
  nand g44 (n_34, n_131, n_132, n_133);
  xor g45 (n_134, A[8], A[4]);
  xor g46 (n_96, n_134, A[1]);
  nand g47 (n_135, A[8], A[4]);
  nand g48 (n_136, A[1], A[4]);
  nand g5 (n_137, A[8], A[1]);
  nand g49 (n_97, n_135, n_136, n_137);
  xor g50 (n_138, A[2], n_95);
  xor g51 (n_59, n_138, n_96);
  nand g52 (n_139, A[2], n_95);
  nand g53 (n_140, n_96, n_95);
  nand g54 (n_141, A[2], n_96);
  nand g6 (n_33, n_139, n_140, n_141);
  xor g55 (n_142, A[9], A[5]);
  xor g56 (n_98, n_142, A[2]);
  nand g57 (n_143, A[9], A[5]);
  nand g58 (n_144, A[2], A[5]);
  nand g59 (n_145, A[9], A[2]);
  nand g60 (n_99, n_143, n_144, n_145);
  xor g61 (n_146, A[3], n_97);
  xor g62 (n_58, n_146, n_98);
  nand g63 (n_147, A[3], n_97);
  nand g64 (n_148, n_98, n_97);
  nand g65 (n_149, A[3], n_98);
  nand g66 (n_32, n_147, n_148, n_149);
  xor g67 (n_150, A[10], A[6]);
  xor g68 (n_100, n_150, A[3]);
  nand g69 (n_151, A[10], A[6]);
  nand g70 (n_152, A[3], A[6]);
  nand g71 (n_153, A[10], A[3]);
  nand g72 (n_101, n_151, n_152, n_153);
  xor g73 (n_154, A[4], n_99);
  xor g74 (n_57, n_154, n_100);
  nand g75 (n_155, A[4], n_99);
  nand g76 (n_156, n_100, n_99);
  nand g77 (n_157, A[4], n_100);
  nand g78 (n_31, n_155, n_156, n_157);
  xor g79 (n_158, A[11], A[7]);
  xor g80 (n_102, n_158, A[4]);
  nand g81 (n_159, A[11], A[7]);
  nand g82 (n_160, A[4], A[7]);
  nand g83 (n_161, A[11], A[4]);
  nand g84 (n_103, n_159, n_160, n_161);
  xor g85 (n_162, A[5], n_101);
  xor g86 (n_56, n_162, n_102);
  nand g87 (n_163, A[5], n_101);
  nand g88 (n_164, n_102, n_101);
  nand g89 (n_165, A[5], n_102);
  nand g90 (n_30, n_163, n_164, n_165);
  xor g91 (n_166, A[12], A[8]);
  xor g92 (n_104, n_166, A[5]);
  nand g93 (n_167, A[12], A[8]);
  nand g94 (n_168, A[5], A[8]);
  nand g95 (n_169, A[12], A[5]);
  nand g96 (n_105, n_167, n_168, n_169);
  xor g97 (n_170, A[6], n_103);
  xor g98 (n_55, n_170, n_104);
  nand g99 (n_171, A[6], n_103);
  nand g100 (n_172, n_104, n_103);
  nand g101 (n_173, A[6], n_104);
  nand g102 (n_29, n_171, n_172, n_173);
  xor g103 (n_174, A[13], A[9]);
  xor g104 (n_106, n_174, A[6]);
  nand g105 (n_175, A[13], A[9]);
  nand g106 (n_176, A[6], A[9]);
  nand g107 (n_177, A[13], A[6]);
  nand g108 (n_107, n_175, n_176, n_177);
  xor g109 (n_178, A[7], n_105);
  xor g110 (n_54, n_178, n_106);
  nand g111 (n_179, A[7], n_105);
  nand g112 (n_180, n_106, n_105);
  nand g113 (n_181, A[7], n_106);
  nand g114 (n_28, n_179, n_180, n_181);
  xor g115 (n_182, A[14], A[10]);
  xor g116 (n_108, n_182, A[7]);
  nand g117 (n_183, A[14], A[10]);
  nand g118 (n_184, A[7], A[10]);
  nand g119 (n_185, A[14], A[7]);
  nand g120 (n_109, n_183, n_184, n_185);
  xor g121 (n_186, A[8], n_107);
  xor g122 (n_53, n_186, n_108);
  nand g123 (n_187, A[8], n_107);
  nand g124 (n_188, n_108, n_107);
  nand g125 (n_189, A[8], n_108);
  nand g126 (n_27, n_187, n_188, n_189);
  xor g127 (n_190, A[15], A[11]);
  xor g128 (n_110, n_190, A[8]);
  nand g129 (n_191, A[15], A[11]);
  nand g130 (n_192, A[8], A[11]);
  nand g131 (n_193, A[15], A[8]);
  nand g132 (n_38, n_191, n_192, n_193);
  xor g133 (n_194, A[9], n_109);
  xor g134 (n_52, n_194, n_110);
  nand g135 (n_195, A[9], n_109);
  nand g136 (n_196, n_110, n_109);
  nand g137 (n_197, A[9], n_110);
  nand g138 (n_26, n_195, n_196, n_197);
  nand g145 (n_201, A[9], A[10]);
  xor g147 (n_202, n_37, n_38);
  xor g148 (n_51, n_202, n_39);
  nand g149 (n_203, n_37, n_38);
  nand g150 (n_204, n_39, n_38);
  nand g151 (n_205, n_37, n_39);
  nand g152 (n_25, n_203, n_204, n_205);
  xor g153 (n_42, A[13], A[11]);
  and g154 (n_114, A[13], A[11]);
  nand g158 (n_208, n_41, A[10]);
  xor g161 (n_210, n_42, n_111);
  xor g162 (n_50, n_210, n_112);
  nand g163 (n_211, n_42, n_111);
  nand g164 (n_212, n_112, n_111);
  nand g165 (n_213, n_42, n_112);
  nand g166 (n_24, n_211, n_212, n_213);
  xor g167 (n_115, A[14], A[12]);
  and g168 (n_119, A[14], A[12]);
  nand g172 (n_216, n_114, A[11]);
  xor g175 (n_218, n_115, n_116);
  xor g176 (n_49, n_218, n_117);
  nand g177 (n_219, n_115, n_116);
  nand g178 (n_220, n_117, n_116);
  nand g179 (n_221, n_115, n_117);
  nand g180 (n_23, n_219, n_220, n_221);
  xor g181 (n_120, A[15], A[13]);
  and g182 (n_123, A[15], A[13]);
  nand g186 (n_224, n_119, A[12]);
  xor g189 (n_226, n_120, n_121);
  xor g190 (n_48, n_226, n_122);
  nand g191 (n_227, n_120, n_121);
  nand g192 (n_228, n_122, n_121);
  nand g193 (n_229, n_120, n_122);
  nand g194 (n_22, n_227, n_228, n_229);
  xor g196 (n_124, n_230, A[13]);
  nand g198 (n_232, A[13], A[14]);
  nand g200 (n_128, n_231, n_232, n_233);
  xor g201 (n_234, n_123, n_124);
  xor g202 (n_47, n_234, n_125);
  nand g203 (n_235, n_123, n_124);
  nand g204 (n_236, n_125, n_124);
  nand g205 (n_237, n_123, n_125);
  nand g206 (n_46, n_235, n_236, n_237);
  xor g207 (n_127, A[15], A[14]);
  and g208 (n_129, A[15], A[14]);
  nand g212 (n_240, n_128, n_127);
  xor g216 (n_20, n_242, n_129);
  nand g218 (n_244, n_129, A[15]);
  nand g220 (n_44, n_243, n_244, n_245);
  nand g28 (n_268, A[4], A[0]);
  xor g32 (Z[4], A[4], A[0]);
  nand g34 (n_273, A[5], A[1]);
  nand g37 (n_277, n_273, n_274, n_275);
  xor g226 (n_276, A[5], A[1]);
  nand g228 (n_278, A[2], n_61);
  nand g229 (n_279, A[2], n_277);
  nand g230 (n_280, n_61, n_277);
  nand g231 (n_282, n_278, n_279, n_280);
  xor g232 (n_281, A[2], n_61);
  xor g233 (Z[6], n_277, n_281);
  nand g234 (n_283, n_35, n_60);
  nand g235 (n_284, n_35, n_282);
  nand g236 (n_285, n_60, n_282);
  nand g237 (n_287, n_283, n_284, n_285);
  xor g238 (n_286, n_35, n_60);
  xor g239 (Z[7], n_282, n_286);
  nand g240 (n_288, n_34, n_59);
  nand g241 (n_289, n_34, n_287);
  nand g242 (n_290, n_59, n_287);
  nand g243 (n_292, n_288, n_289, n_290);
  xor g244 (n_291, n_34, n_59);
  xor g245 (Z[8], n_287, n_291);
  nand g246 (n_293, n_33, n_58);
  nand g247 (n_294, n_33, n_292);
  nand g248 (n_295, n_58, n_292);
  nand g249 (n_297, n_293, n_294, n_295);
  xor g250 (n_296, n_33, n_58);
  xor g251 (Z[9], n_292, n_296);
  nand g252 (n_298, n_32, n_57);
  nand g253 (n_299, n_32, n_297);
  nand g254 (n_300, n_57, n_297);
  nand g255 (n_302, n_298, n_299, n_300);
  xor g256 (n_301, n_32, n_57);
  xor g257 (Z[10], n_297, n_301);
  nand g258 (n_303, n_31, n_56);
  nand g259 (n_304, n_31, n_302);
  nand g260 (n_305, n_56, n_302);
  nand g261 (n_307, n_303, n_304, n_305);
  xor g262 (n_306, n_31, n_56);
  xor g263 (Z[11], n_302, n_306);
  nand g264 (n_308, n_30, n_55);
  nand g265 (n_309, n_30, n_307);
  nand g266 (n_310, n_55, n_307);
  nand g267 (n_312, n_308, n_309, n_310);
  xor g268 (n_311, n_30, n_55);
  xor g269 (Z[12], n_307, n_311);
  nand g270 (n_313, n_29, n_54);
  nand g271 (n_314, n_29, n_312);
  nand g272 (n_315, n_54, n_312);
  nand g273 (n_317, n_313, n_314, n_315);
  xor g274 (n_316, n_29, n_54);
  xor g275 (Z[13], n_312, n_316);
  nand g276 (n_318, n_28, n_53);
  nand g277 (n_319, n_28, n_317);
  nand g278 (n_320, n_53, n_317);
  nand g279 (n_322, n_318, n_319, n_320);
  xor g280 (n_321, n_28, n_53);
  xor g281 (Z[14], n_317, n_321);
  nand g282 (n_323, n_27, n_52);
  nand g283 (n_324, n_27, n_322);
  nand g284 (n_325, n_52, n_322);
  nand g285 (n_327, n_323, n_324, n_325);
  xor g286 (n_326, n_27, n_52);
  xor g287 (Z[15], n_322, n_326);
  nand g288 (n_328, n_26, n_51);
  nand g289 (n_329, n_26, n_327);
  nand g290 (n_330, n_51, n_327);
  nand g291 (n_332, n_328, n_329, n_330);
  xor g292 (n_331, n_26, n_51);
  xor g293 (Z[16], n_327, n_331);
  nand g294 (n_333, n_25, n_50);
  nand g295 (n_334, n_25, n_332);
  nand g296 (n_335, n_50, n_332);
  nand g297 (n_337, n_333, n_334, n_335);
  xor g298 (n_336, n_25, n_50);
  xor g299 (Z[17], n_332, n_336);
  nand g300 (n_338, n_24, n_49);
  nand g301 (n_339, n_24, n_337);
  nand g302 (n_340, n_49, n_337);
  nand g303 (n_342, n_338, n_339, n_340);
  xor g304 (n_341, n_24, n_49);
  xor g305 (Z[18], n_337, n_341);
  nand g306 (n_343, n_23, n_48);
  nand g307 (n_344, n_23, n_342);
  nand g308 (n_345, n_48, n_342);
  nand g309 (n_347, n_343, n_344, n_345);
  xor g310 (n_346, n_23, n_48);
  xor g311 (Z[19], n_342, n_346);
  nand g312 (n_348, n_22, n_47);
  nand g313 (n_349, n_22, n_347);
  nand g314 (n_350, n_47, n_347);
  nand g315 (n_352, n_348, n_349, n_350);
  xor g316 (n_351, n_22, n_47);
  xor g317 (Z[20], n_347, n_351);
  nand g318 (n_353, n_21, n_46);
  nand g319 (n_354, n_21, n_352);
  nand g320 (n_355, n_46, n_352);
  nand g321 (n_357, n_353, n_354, n_355);
  xor g322 (n_356, n_21, n_46);
  xor g323 (Z[21], n_352, n_356);
  nand g324 (n_358, n_20, n_45);
  nand g325 (n_359, n_20, n_357);
  nand g326 (n_360, n_45, n_357);
  nand g327 (n_362, n_358, n_359, n_360);
  xor g328 (n_361, n_20, n_45);
  xor g329 (Z[22], n_357, n_361);
  nand g332 (n_365, n_44, n_362);
  nand g333 (n_367, n_363, n_364, n_365);
  xor g335 (Z[23], n_362, n_366);
  xnor g342 (n_37, A[16], A[12]);
  and g343 (n_41, A[12], wc);
  not gc (wc, A[16]);
  xnor g344 (n_39, A[10], A[9]);
  or g345 (n_111, A[9], A[10], wc0);
  not gc0 (wc0, n_201);
  xnor g346 (n_116, n_114, A[11]);
  xnor g348 (n_121, n_119, A[12]);
  xnor g350 (n_230, A[16], A[14]);
  or g351 (n_231, wc1, A[16]);
  not gc1 (wc1, A[14]);
  or g352 (n_233, wc2, A[16]);
  not gc2 (wc2, A[13]);
  xnor g354 (n_242, A[16], A[15]);
  or g355 (n_243, wc3, A[16]);
  not gc3 (wc3, A[15]);
  or g356 (n_245, A[16], wc4);
  not gc4 (wc4, n_129);
  xnor g357 (n_112, n_41, A[10]);
  or g359 (n_122, A[11], wc5, n_114);
  not gc5 (wc5, n_216);
  or g360 (n_125, A[12], wc6, n_119);
  not gc6 (wc6, n_224);
  or g361 (n_117, A[10], n_41, wc7);
  not gc7 (wc7, n_208);
  xnor g362 (n_21, n_128, n_127);
  or g364 (n_363, A[16], wc8);
  not gc8 (wc8, n_44);
  xnor g365 (n_366, n_44, A[16]);
  or g366 (n_45, wc9, n_127, n_128);
  not gc9 (wc9, n_240);
  or g368 (n_274, wc10, n_268);
  not gc10 (wc10, A[5]);
  or g369 (n_275, wc11, n_268);
  not gc11 (wc11, A[1]);
  xnor g370 (Z[5], n_268, n_276);
  or g371 (n_364, A[16], wc12);
  not gc12 (wc12, n_362);
  not g372 (Z[24], n_367);
endmodule

module mult_signed_const_107_GENERIC(A, Z);
  input [16:0] A;
  output [24:0] Z;
  wire [16:0] A;
  wire [24:0] Z;
  mult_signed_const_107_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_175_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * -1899;"
  input [16:0] A;
  output [28:0] Z;
  wire [16:0] A;
  wire [28:0] Z;
  wire n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_39, n_40, n_41, n_42, n_43, n_46, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_110, n_112, n_113;
  wire n_115, n_116, n_118, n_119, n_121, n_122, n_123, n_125;
  wire n_126, n_127, n_128, n_130, n_131, n_132, n_134, n_135;
  wire n_136, n_137, n_140, n_141, n_143, n_144, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_190, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_201, n_202, n_203;
  wire n_204, n_206, n_208, n_210, n_211, n_212, n_218, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_306, n_307;
  wire n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_335, n_336, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_367;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_381, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_422, n_424, n_425, n_426;
  wire n_427, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_438, n_440, n_441, n_442, n_443, n_451, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567;
  wire n_568, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_580, n_582, n_583, n_585;
  assign Z[0] = A[0];
  xor g94 (n_72, A[0], n_110);
  xor g102 (n_71, n_220, n_113);
  nand g104 (n_222, n_113, n_112);
  nand g106 (n_41, n_221, n_222, n_223);
  xor g108 (n_116, n_224, A[0]);
  nand g112 (n_118, n_225, n_226, n_227);
  xor g114 (n_70, n_228, n_116);
  nand g116 (n_230, n_116, n_115);
  nand g118 (n_40, n_229, n_230, n_231);
  xor g120 (n_119, n_232, A[1]);
  nand g124 (n_122, n_233, n_234, n_235);
  xor g126 (n_69, n_236, n_119);
  nand g128 (n_238, n_119, n_118);
  nand g130 (n_39, n_237, n_238, n_239);
  xor g133 (n_240, A[2], A[0]);
  nand g135 (n_241, A[2], A[0]);
  nand g138 (n_126, n_241, n_226, n_243);
  xor g139 (n_244, n_121, n_122);
  xor g140 (n_68, n_244, n_123);
  nand g141 (n_245, n_121, n_122);
  nand g142 (n_246, n_123, n_122);
  nand g143 (n_247, n_121, n_123);
  nand g144 (n_38, n_245, n_246, n_247);
  xor g146 (n_127, n_248, A[3]);
  nand g150 (n_130, n_249, n_250, n_251);
  xor g152 (n_128, n_252, n_125);
  nand g155 (n_255, A[1], n_125);
  nand g156 (n_46, n_234, n_254, n_255);
  xor g157 (n_256, n_126, n_127);
  xor g158 (n_67, n_256, n_128);
  nand g159 (n_257, n_126, n_127);
  nand g160 (n_258, n_128, n_127);
  nand g161 (n_259, n_126, n_128);
  nand g162 (n_37, n_257, n_258, n_259);
  xor g164 (n_131, n_260, A[4]);
  nand g168 (n_134, n_261, n_262, n_263);
  xor g170 (n_132, n_264, n_130);
  nand g173 (n_267, A[2], n_130);
  nand g174 (n_137, n_265, n_266, n_267);
  xor g175 (n_268, n_131, n_46);
  xor g176 (n_66, n_268, n_132);
  nand g177 (n_269, n_131, n_46);
  nand g178 (n_270, n_132, n_46);
  nand g179 (n_271, n_131, n_132);
  nand g180 (n_36, n_269, n_270, n_271);
  xor g182 (n_135, n_272, A[5]);
  nand g186 (n_140, n_273, n_274, n_275);
  xor g188 (n_136, n_276, n_134);
  nand g191 (n_279, A[3], n_134);
  nand g192 (n_143, n_250, n_278, n_279);
  xor g193 (n_280, n_135, n_136);
  xor g194 (n_65, n_280, n_137);
  nand g195 (n_281, n_135, n_136);
  nand g196 (n_282, n_137, n_136);
  nand g197 (n_283, n_135, n_137);
  nand g198 (n_35, n_281, n_282, n_283);
  xor g200 (n_141, n_284, A[6]);
  nand g204 (n_147, n_285, n_286, n_287);
  xor g212 (n_144, n_292, n_141);
  nand g214 (n_294, n_141, n_140);
  nand g216 (n_151, n_293, n_294, n_295);
  xor g218 (n_64, n_296, n_144);
  nand g220 (n_298, n_144, n_143);
  nand g222 (n_34, n_297, n_298, n_299);
  xor g224 (n_148, n_300, A[7]);
  nand g228 (n_154, n_301, n_302, n_303);
  nand g234 (n_153, n_274, n_306, n_307);
  xor g235 (n_308, n_146, n_147);
  xor g236 (n_150, n_308, n_148);
  nand g237 (n_309, n_146, n_147);
  nand g238 (n_310, n_148, n_147);
  nand g239 (n_311, n_146, n_148);
  nand g240 (n_158, n_309, n_310, n_311);
  xor g241 (n_312, n_149, n_150);
  xor g242 (n_63, n_312, n_151);
  nand g243 (n_313, n_149, n_150);
  nand g244 (n_314, n_151, n_150);
  nand g245 (n_315, n_149, n_151);
  nand g246 (n_33, n_313, n_314, n_315);
  xor g248 (n_155, n_316, A[8]);
  nand g252 (n_161, n_317, n_318, n_319);
  nand g258 (n_160, n_286, n_322, n_323);
  xor g259 (n_324, n_153, n_154);
  xor g260 (n_157, n_324, n_155);
  nand g261 (n_325, n_153, n_154);
  nand g262 (n_326, n_155, n_154);
  nand g263 (n_327, n_153, n_155);
  nand g264 (n_165, n_325, n_326, n_327);
  xor g265 (n_328, n_156, n_157);
  xor g266 (n_62, n_328, n_158);
  nand g267 (n_329, n_156, n_157);
  nand g268 (n_330, n_158, n_157);
  nand g269 (n_331, n_156, n_158);
  nand g270 (n_32, n_329, n_330, n_331);
  xor g272 (n_162, n_332, A[9]);
  nand g276 (n_168, n_333, n_334, n_335);
  nand g282 (n_167, n_302, n_338, n_339);
  xor g283 (n_340, n_160, n_161);
  xor g284 (n_164, n_340, n_162);
  nand g285 (n_341, n_160, n_161);
  nand g286 (n_342, n_162, n_161);
  nand g287 (n_343, n_160, n_162);
  nand g288 (n_172, n_341, n_342, n_343);
  xor g289 (n_344, n_163, n_164);
  xor g290 (n_61, n_344, n_165);
  nand g291 (n_345, n_163, n_164);
  nand g292 (n_346, n_165, n_164);
  nand g293 (n_347, n_163, n_165);
  nand g294 (n_31, n_345, n_346, n_347);
  xor g296 (n_169, n_348, A[10]);
  nand g300 (n_175, n_349, n_350, n_351);
  nand g306 (n_176, n_318, n_354, n_355);
  xor g307 (n_356, n_167, n_168);
  xor g308 (n_171, n_356, n_169);
  nand g309 (n_357, n_167, n_168);
  nand g310 (n_358, n_169, n_168);
  nand g311 (n_359, n_167, n_169);
  nand g312 (n_180, n_357, n_358, n_359);
  xor g313 (n_360, n_170, n_171);
  xor g314 (n_60, n_360, n_172);
  nand g315 (n_361, n_170, n_171);
  nand g316 (n_362, n_172, n_171);
  nand g317 (n_363, n_170, n_172);
  nand g318 (n_30, n_361, n_362, n_363);
  xor g321 (n_364, A[11], A[9]);
  nand g323 (n_365, A[11], A[9]);
  nand g326 (n_182, n_365, n_334, n_367);
  xor g328 (n_178, A[5], n_174);
  xor g333 (n_372, n_175, n_176);
  xor g334 (n_179, n_372, n_177);
  nand g335 (n_373, n_175, n_176);
  nand g336 (n_374, n_177, n_176);
  nand g337 (n_375, n_175, n_177);
  nand g338 (n_186, n_373, n_374, n_375);
  xor g339 (n_376, n_178, n_179);
  xor g340 (n_59, n_376, n_180);
  nand g341 (n_377, n_178, n_179);
  nand g342 (n_378, n_180, n_179);
  nand g343 (n_379, n_178, n_180);
  nand g344 (n_29, n_377, n_378, n_379);
  nand g349 (n_383, A[16], A[10]);
  nand g350 (n_190, n_381, n_350, n_383);
  xor g352 (n_185, n_384, n_181);
  nand g354 (n_386, n_181, A[12]);
  nand g356 (n_192, n_385, n_386, n_387);
  xor g357 (n_388, n_182, n_183);
  xor g358 (n_187, n_388, n_184);
  nand g359 (n_389, n_182, n_183);
  nand g360 (n_390, n_184, n_183);
  nand g361 (n_391, n_182, n_184);
  nand g362 (n_194, n_389, n_390, n_391);
  xor g363 (n_392, n_185, n_186);
  xor g364 (n_58, n_392, n_187);
  nand g365 (n_393, n_185, n_186);
  nand g366 (n_394, n_187, n_186);
  nand g367 (n_395, n_185, n_187);
  nand g368 (n_28, n_393, n_394, n_395);
  nand g382 (n_199, n_401, n_402, n_403);
  xor g383 (n_404, n_192, n_193);
  xor g384 (n_57, n_404, n_194);
  nand g385 (n_405, n_192, n_193);
  nand g386 (n_406, n_194, n_193);
  nand g387 (n_407, n_192, n_194);
  nand g388 (n_56, n_405, n_406, n_407);
  xor g389 (n_408, A[16], A[14]);
  nand g391 (n_409, A[16], A[14]);
  nand g394 (n_202, n_409, n_410, n_411);
  xor g395 (n_412, A[12], n_195);
  xor g396 (n_198, n_412, n_196);
  nand g397 (n_413, A[12], n_195);
  nand g398 (n_414, n_196, n_195);
  nand g399 (n_415, A[12], n_196);
  nand g400 (n_204, n_413, n_414, n_415);
  xor g401 (n_416, n_197, n_198);
  xor g402 (n_27, n_416, n_199);
  nand g403 (n_417, n_197, n_198);
  nand g404 (n_418, n_199, n_198);
  nand g405 (n_419, n_197, n_199);
  nand g406 (n_55, n_417, n_418, n_419);
  xor g407 (n_201, A[15], A[13]);
  and g408 (n_206, A[15], A[13]);
  xor g410 (n_203, A[9], n_201);
  xor g415 (n_424, n_202, n_203);
  xor g416 (n_26, n_424, n_204);
  nand g417 (n_425, n_202, n_203);
  nand g418 (n_426, n_204, n_203);
  nand g419 (n_427, n_202, n_204);
  nand g420 (n_54, n_425, n_426, n_427);
  nand g426 (n_211, n_429, n_430, n_431);
  xor g428 (n_25, n_432, n_208);
  nand g431 (n_435, n_206, n_208);
  nand g432 (n_53, n_433, n_434, n_435);
  nand g438 (n_438, n_211, n_210);
  xor g442 (n_23, n_440, n_212);
  nand g446 (n_51, n_441, n_442, n_443);
  nand g18 (n_458, n_73, n_455);
  nand g19 (n_460, n_456, n_457, n_458);
  xor g21 (Z[2], n_455, n_459);
  nand g22 (n_461, n_43, n_72);
  nand g23 (n_462, n_43, n_460);
  nand g24 (n_463, n_72, n_460);
  nand g25 (n_465, n_461, n_462, n_463);
  xor g26 (n_464, n_43, n_72);
  xor g27 (Z[3], n_460, n_464);
  nand g28 (n_466, n_42, n_71);
  nand g29 (n_467, n_42, n_465);
  nand g30 (n_468, n_71, n_465);
  nand g31 (n_470, n_466, n_467, n_468);
  xor g32 (n_469, n_42, n_71);
  xor g33 (Z[4], n_465, n_469);
  nand g34 (n_471, n_41, n_70);
  nand g35 (n_472, n_41, n_470);
  nand g36 (n_473, n_70, n_470);
  nand g37 (n_475, n_471, n_472, n_473);
  xor g38 (n_474, n_41, n_70);
  xor g39 (Z[5], n_470, n_474);
  nand g40 (n_476, n_40, n_69);
  nand g41 (n_477, n_40, n_475);
  nand g42 (n_478, n_69, n_475);
  nand g43 (n_480, n_476, n_477, n_478);
  xor g44 (n_479, n_40, n_69);
  xor g45 (Z[6], n_475, n_479);
  nand g46 (n_481, n_39, n_68);
  nand g47 (n_482, n_39, n_480);
  nand g48 (n_483, n_68, n_480);
  nand g49 (n_485, n_481, n_482, n_483);
  xor g50 (n_484, n_39, n_68);
  xor g51 (Z[7], n_480, n_484);
  nand g52 (n_486, n_38, n_67);
  nand g53 (n_487, n_38, n_485);
  nand g54 (n_488, n_67, n_485);
  nand g55 (n_490, n_486, n_487, n_488);
  xor g56 (n_489, n_38, n_67);
  xor g57 (Z[8], n_485, n_489);
  nand g58 (n_491, n_37, n_66);
  nand g59 (n_492, n_37, n_490);
  nand g60 (n_493, n_66, n_490);
  nand g61 (n_495, n_491, n_492, n_493);
  xor g62 (n_494, n_37, n_66);
  xor g63 (Z[9], n_490, n_494);
  nand g64 (n_496, n_36, n_65);
  nand g65 (n_497, n_36, n_495);
  nand g66 (n_498, n_65, n_495);
  nand g67 (n_500, n_496, n_497, n_498);
  xor g68 (n_499, n_36, n_65);
  xor g69 (Z[10], n_495, n_499);
  nand g70 (n_501, n_35, n_64);
  nand g71 (n_502, n_35, n_500);
  nand g72 (n_503, n_64, n_500);
  nand g73 (n_505, n_501, n_502, n_503);
  xor g74 (n_504, n_35, n_64);
  xor g75 (Z[11], n_500, n_504);
  nand g76 (n_506, n_34, n_63);
  nand g77 (n_507, n_34, n_505);
  nand g78 (n_508, n_63, n_505);
  nand g79 (n_510, n_506, n_507, n_508);
  xor g80 (n_509, n_34, n_63);
  xor g81 (Z[12], n_505, n_509);
  nand g82 (n_511, n_33, n_62);
  nand g83 (n_512, n_33, n_510);
  nand g84 (n_513, n_62, n_510);
  nand g85 (n_515, n_511, n_512, n_513);
  xor g86 (n_514, n_33, n_62);
  xor g469 (Z[13], n_510, n_514);
  nand g470 (n_516, n_32, n_61);
  nand g471 (n_517, n_32, n_515);
  nand g472 (n_518, n_61, n_515);
  nand g473 (n_520, n_516, n_517, n_518);
  xor g474 (n_519, n_32, n_61);
  xor g475 (Z[14], n_515, n_519);
  nand g476 (n_521, n_31, n_60);
  nand g477 (n_522, n_31, n_520);
  nand g478 (n_523, n_60, n_520);
  nand g479 (n_525, n_521, n_522, n_523);
  xor g480 (n_524, n_31, n_60);
  xor g481 (Z[15], n_520, n_524);
  nand g482 (n_526, n_30, n_59);
  nand g483 (n_527, n_30, n_525);
  nand g484 (n_528, n_59, n_525);
  nand g485 (n_530, n_526, n_527, n_528);
  xor g486 (n_529, n_30, n_59);
  xor g487 (Z[16], n_525, n_529);
  nand g488 (n_531, n_29, n_58);
  nand g489 (n_532, n_29, n_530);
  nand g490 (n_533, n_58, n_530);
  nand g491 (n_535, n_531, n_532, n_533);
  xor g492 (n_534, n_29, n_58);
  xor g493 (Z[17], n_530, n_534);
  nand g494 (n_536, n_28, n_57);
  nand g495 (n_537, n_28, n_535);
  nand g496 (n_538, n_57, n_535);
  nand g497 (n_540, n_536, n_537, n_538);
  xor g498 (n_539, n_28, n_57);
  xor g499 (Z[18], n_535, n_539);
  nand g500 (n_541, n_27, n_56);
  nand g501 (n_542, n_27, n_540);
  nand g502 (n_543, n_56, n_540);
  nand g503 (n_545, n_541, n_542, n_543);
  xor g504 (n_544, n_27, n_56);
  xor g505 (Z[19], n_540, n_544);
  nand g506 (n_546, n_26, n_55);
  nand g507 (n_547, n_26, n_545);
  nand g508 (n_548, n_55, n_545);
  nand g509 (n_550, n_546, n_547, n_548);
  xor g510 (n_549, n_26, n_55);
  xor g511 (Z[20], n_545, n_549);
  nand g512 (n_551, n_25, n_54);
  nand g513 (n_552, n_25, n_550);
  nand g514 (n_553, n_54, n_550);
  nand g515 (n_555, n_551, n_552, n_553);
  xor g516 (n_554, n_25, n_54);
  xor g517 (Z[21], n_550, n_554);
  nand g518 (n_556, n_24, n_53);
  nand g519 (n_557, n_24, n_555);
  nand g520 (n_558, n_53, n_555);
  nand g521 (n_560, n_556, n_557, n_558);
  xor g522 (n_559, n_24, n_53);
  xor g523 (Z[22], n_555, n_559);
  nand g524 (n_561, n_23, n_52);
  nand g525 (n_562, n_23, n_560);
  nand g526 (n_563, n_52, n_560);
  nand g527 (n_565, n_561, n_562, n_563);
  xor g528 (n_564, n_23, n_52);
  xor g529 (Z[23], n_560, n_564);
  nand g530 (n_566, A[13], n_51);
  nand g531 (n_567, A[13], n_565);
  nand g532 (n_568, n_51, n_565);
  nand g533 (n_570, n_566, n_567, n_568);
  xor g534 (n_569, A[13], n_51);
  xor g535 (Z[24], n_565, n_569);
  nand g538 (n_573, A[14], n_570);
  nand g539 (n_575, n_571, n_572, n_573);
  nand g544 (n_578, A[15], n_575);
  nand g545 (n_580, n_576, n_577, n_578);
  nand g549 (n_582, A[16], n_580);
  xor g553 (Z[27], n_580, n_174);
  xor g556 (n_73, A[2], A[1]);
  nor g557 (n_43, A[2], A[1]);
  xor g558 (n_110, A[3], A[2]);
  nor g559 (n_113, A[3], A[2]);
  xor g560 (n_112, A[4], A[3]);
  nor g561 (n_115, A[4], A[3]);
  xor g562 (n_224, A[5], A[4]);
  or g563 (n_225, A[5], A[4]);
  or g564 (n_226, wc, A[4]);
  not gc (wc, A[0]);
  or g565 (n_227, wc0, A[5]);
  not gc0 (wc0, A[0]);
  xor g566 (n_232, A[6], A[5]);
  or g567 (n_233, A[6], A[5]);
  or g568 (n_234, wc1, A[5]);
  not gc1 (wc1, A[1]);
  or g569 (n_235, wc2, A[6]);
  not gc2 (wc2, A[1]);
  xor g570 (n_121, A[7], A[6]);
  nor g571 (n_125, A[7], A[6]);
  xnor g572 (n_123, n_240, A[4]);
  or g573 (n_243, wc3, A[4]);
  not gc3 (wc3, A[2]);
  xor g574 (n_248, A[8], A[7]);
  or g575 (n_249, A[8], A[7]);
  or g576 (n_250, wc4, A[7]);
  not gc4 (wc4, A[3]);
  or g577 (n_251, wc5, A[8]);
  not gc5 (wc5, A[3]);
  xnor g578 (n_252, A[5], A[1]);
  xor g579 (n_260, A[9], A[8]);
  or g580 (n_261, A[9], A[8]);
  or g581 (n_262, wc6, A[8]);
  not gc6 (wc6, A[4]);
  or g582 (n_263, wc7, A[9]);
  not gc7 (wc7, A[4]);
  xnor g583 (n_264, A[6], A[2]);
  or g584 (n_265, wc8, A[6]);
  not gc8 (wc8, A[2]);
  xor g585 (n_272, A[10], A[9]);
  or g586 (n_273, A[10], A[9]);
  or g587 (n_274, wc9, A[9]);
  not gc9 (wc9, A[5]);
  or g588 (n_275, wc10, A[10]);
  not gc10 (wc10, A[5]);
  xnor g589 (n_276, A[7], A[3]);
  xor g590 (n_284, A[11], A[10]);
  or g591 (n_285, A[11], A[10]);
  or g592 (n_286, wc11, A[10]);
  not gc11 (wc11, A[6]);
  or g593 (n_287, wc12, A[11]);
  not gc12 (wc12, A[6]);
  xnor g594 (n_288, A[8], A[4]);
  xor g595 (n_300, A[12], A[11]);
  or g596 (n_301, A[12], A[11]);
  or g597 (n_302, wc13, A[11]);
  not gc13 (wc13, A[7]);
  or g598 (n_303, wc14, A[12]);
  not gc14 (wc14, A[7]);
  xnor g599 (n_304, A[9], A[5]);
  or g600 (n_306, A[9], A[1]);
  or g601 (n_307, A[1], wc15);
  not gc15 (wc15, A[5]);
  xor g602 (n_316, A[13], A[12]);
  or g603 (n_317, A[13], A[12]);
  or g604 (n_318, wc16, A[12]);
  not gc16 (wc16, A[8]);
  or g605 (n_319, wc17, A[13]);
  not gc17 (wc17, A[8]);
  xnor g606 (n_320, A[10], A[6]);
  or g607 (n_322, A[10], A[2]);
  or g608 (n_323, A[2], wc18);
  not gc18 (wc18, A[6]);
  xor g609 (n_332, A[14], A[13]);
  or g610 (n_333, A[14], A[13]);
  or g611 (n_334, wc19, A[13]);
  not gc19 (wc19, A[9]);
  or g612 (n_335, wc20, A[14]);
  not gc20 (wc20, A[9]);
  xnor g613 (n_336, A[11], A[7]);
  or g614 (n_338, A[11], A[3]);
  or g615 (n_339, A[3], wc21);
  not gc21 (wc21, A[7]);
  xor g616 (n_348, A[15], A[14]);
  or g617 (n_349, A[15], A[14]);
  or g618 (n_350, wc22, A[14]);
  not gc22 (wc22, A[10]);
  or g619 (n_351, wc23, A[15]);
  not gc23 (wc23, A[10]);
  xnor g620 (n_352, A[12], A[8]);
  or g621 (n_354, A[12], A[4]);
  or g622 (n_355, A[4], wc24);
  not gc24 (wc24, A[8]);
  xnor g623 (n_174, A[16], A[15]);
  and g624 (n_181, wc25, A[16]);
  not gc25 (wc25, A[15]);
  xnor g625 (n_177, n_364, A[13]);
  or g626 (n_367, wc26, A[13]);
  not gc26 (wc26, A[11]);
  or g628 (n_381, A[14], wc27);
  not gc27 (wc27, A[16]);
  xnor g629 (n_384, A[12], A[6]);
  or g630 (n_385, A[6], wc28);
  not gc28 (wc28, A[12]);
  and g632 (n_195, A[13], wc29);
  not gc29 (wc29, A[15]);
  or g633 (n_399, A[7], wc30);
  not gc30 (wc30, A[11]);
  xnor g634 (n_197, n_408, A[8]);
  or g635 (n_410, A[8], wc31);
  not gc31 (wc31, A[14]);
  or g636 (n_411, A[8], wc32);
  not gc32 (wc32, A[16]);
  or g637 (n_422, A[9], wc33);
  not gc33 (wc33, n_201);
  or g638 (n_429, wc34, A[16]);
  not gc34 (wc34, A[14]);
  or g639 (n_430, A[10], wc35);
  not gc35 (wc35, A[14]);
  or g640 (n_431, A[16], A[10]);
  xnor g641 (n_210, A[15], A[11]);
  and g642 (n_212, wc36, A[15]);
  not gc36 (wc36, A[11]);
  xor g643 (n_440, A[16], A[12]);
  or g644 (n_441, A[16], A[12]);
  or g645 (n_218, A[0], wc37);
  not gc37 (wc37, n_110);
  xnor g647 (n_220, n_112, A[1]);
  or g648 (n_221, A[1], wc38);
  not gc38 (wc38, n_112);
  or g649 (n_223, A[1], wc39);
  not gc39 (wc39, n_113);
  xnor g650 (n_228, n_115, A[2]);
  or g651 (n_229, A[2], wc40);
  not gc40 (wc40, n_115);
  or g652 (n_254, A[5], wc41);
  not gc41 (wc41, n_125);
  or g654 (n_146, A[4], wc42, wc43);
  not gc43 (wc43, n_262);
  not gc42 (wc42, A[8]);
  xnor g655 (n_149, n_304, A[1]);
  xnor g656 (n_156, n_320, A[2]);
  xnor g657 (n_163, n_336, A[3]);
  xnor g658 (n_170, n_352, A[4]);
  or g660 (n_371, A[5], wc44);
  not gc44 (wc44, n_174);
  xnor g661 (n_183, n_408, A[10]);
  or g662 (n_387, A[6], wc45);
  not gc45 (wc45, n_181);
  or g664 (n_196, wc46, A[11], wc47);
  not gc47 (wc47, n_399);
  not gc46 (wc46, A[7]);
  or g665 (n_208, wc48, wc49, n_201);
  not gc49 (wc49, n_422);
  not gc48 (wc48, A[9]);
  or g668 (n_442, A[12], wc50);
  not gc50 (wc50, n_212);
  or g669 (n_443, A[16], wc51);
  not gc51 (wc51, n_212);
  or g670 (n_451, A[0], wc52);
  not gc52 (wc52, A[1]);
  xnor g671 (n_454, A[1], A[0]);
  or g672 (n_456, A[1], wc53);
  not gc53 (wc53, n_73);
  xnor g673 (n_459, n_73, A[1]);
  or g674 (n_571, A[13], wc54);
  not gc54 (wc54, A[14]);
  or g676 (n_576, A[14], wc55);
  not gc55 (wc55, A[15]);
  or g679 (n_42, wc56, wc57, n_110);
  not gc57 (wc57, n_218);
  not gc56 (wc56, A[0]);
  or g680 (n_231, A[2], wc58);
  not gc58 (wc58, n_116);
  xnor g681 (n_236, n_118, A[3]);
  or g682 (n_237, A[3], wc59);
  not gc59 (wc59, n_118);
  or g683 (n_239, A[3], wc60);
  not gc60 (wc60, n_119);
  or g684 (n_266, A[6], wc61);
  not gc61 (wc61, n_130);
  or g685 (n_278, A[7], wc62);
  not gc62 (wc62, n_134);
  xnor g686 (n_292, n_140, A[0]);
  or g687 (n_293, A[0], wc63);
  not gc63 (wc63, n_140);
  or g688 (n_295, A[0], wc64);
  not gc64 (wc64, n_141);
  or g689 (n_184, wc65, wc66, n_174);
  not gc66 (wc66, n_371);
  not gc65 (wc65, A[5]);
  xnor g690 (n_400, n_190, n_201);
  or g691 (n_401, n_201, wc67);
  not gc67 (wc67, n_190);
  or g692 (n_402, n_336, wc68);
  not gc68 (wc68, n_190);
  or g693 (n_403, n_201, n_336);
  xnor g694 (n_432, n_206, n_183);
  or g695 (n_433, n_183, wc69);
  not gc69 (wc69, n_206);
  or g696 (n_434, wc70, n_183);
  not gc70 (wc70, n_208);
  xnor g697 (n_24, n_211, n_210);
  xnor g699 (Z[1], n_454, A[0]);
  xnor g700 (n_193, n_336, n_400);
  or g701 (n_52, n_210, wc71, n_211);
  not gc71 (wc71, n_438);
  nand g702 (n_455, n_451, A[0]);
  xnor g703 (n_296, n_143, n_288);
  or g704 (n_297, n_288, wc72);
  not gc72 (wc72, n_143);
  or g705 (n_299, n_288, wc73);
  not gc73 (wc73, n_144);
  or g706 (n_457, A[1], wc74);
  not gc74 (wc74, n_455);
  or g707 (n_572, A[13], wc75);
  not gc75 (wc75, n_570);
  xnor g708 (Z[25], n_570, n_332);
  or g709 (n_577, A[14], wc76);
  not gc76 (wc76, n_575);
  xnor g710 (Z[26], n_575, n_348);
  or g711 (n_583, A[15], wc77);
  not gc77 (wc77, n_580);
  or g712 (n_585, wc78, n_181, wc79);
  not gc79 (wc79, n_582);
  not gc78 (wc78, n_583);
  not g713 (Z[28], n_585);
endmodule

module mult_signed_const_175_GENERIC(A, Z);
  input [16:0] A;
  output [28:0] Z;
  wire [16:0] A;
  wire [28:0] Z;
  mult_signed_const_175_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_241_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 1449;"
  input [16:0] A;
  output [27:0] Z;
  wire [16:0] A;
  wire [27:0] Z;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_41, n_42, n_43, n_44, n_45;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_120, n_121;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_174;
  wire n_175, n_176, n_177, n_178, n_180, n_182, n_183, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203;
  wire n_204, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_272, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_317, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_333, n_336;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_349, n_352, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_365, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_404, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_414, n_415, n_416, n_417, n_420, n_421, n_445;
  wire n_446, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_555, n_556, n_558;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  assign Z[2] = A[2];
  xor g69 (n_68, A[5], A[0]);
  and g2 (n_39, A[5], A[0]);
  xor g70 (n_194, A[6], A[3]);
  xor g71 (n_67, n_194, A[1]);
  nand g3 (n_195, A[6], A[3]);
  nand g72 (n_196, A[1], A[3]);
  nand g73 (n_197, A[6], A[1]);
  nand g74 (n_38, n_195, n_196, n_197);
  xor g75 (n_103, A[7], A[4]);
  and g76 (n_105, A[7], A[4]);
  xor g77 (n_198, A[0], A[2]);
  xor g78 (n_66, n_198, n_103);
  nand g79 (n_199, A[0], A[2]);
  nand g4 (n_200, n_103, A[2]);
  nand g5 (n_201, A[0], n_103);
  nand g80 (n_37, n_199, n_200, n_201);
  xor g81 (n_104, A[8], A[5]);
  and g82 (n_107, A[8], A[5]);
  xor g83 (n_202, A[1], A[0]);
  xor g84 (n_106, n_202, A[3]);
  nand g85 (n_203, A[1], A[0]);
  nand g86 (n_204, A[3], A[0]);
  nand g6 (n_108, n_203, n_204, n_196);
  xor g88 (n_206, n_104, n_105);
  xor g89 (n_65, n_206, n_106);
  nand g90 (n_207, n_104, n_105);
  nand g91 (n_208, n_106, n_105);
  nand g92 (n_209, n_104, n_106);
  nand g93 (n_36, n_207, n_208, n_209);
  xor g94 (n_210, A[9], A[6]);
  xor g95 (n_109, n_210, A[2]);
  nand g96 (n_211, A[9], A[6]);
  nand g97 (n_212, A[2], A[6]);
  nand g98 (n_213, A[9], A[2]);
  nand g99 (n_112, n_211, n_212, n_213);
  xor g100 (n_214, A[1], A[4]);
  xor g101 (n_110, n_214, n_107);
  nand g102 (n_215, A[1], A[4]);
  nand g103 (n_216, n_107, A[4]);
  nand g104 (n_217, A[1], n_107);
  nand g105 (n_114, n_215, n_216, n_217);
  xor g106 (n_218, n_108, n_109);
  xor g107 (n_64, n_218, n_110);
  nand g108 (n_219, n_108, n_109);
  nand g109 (n_220, n_110, n_109);
  nand g110 (n_221, n_108, n_110);
  nand g111 (n_35, n_219, n_220, n_221);
  xor g112 (n_111, A[10], A[7]);
  and g113 (n_116, A[10], A[7]);
  xor g114 (n_222, A[3], A[2]);
  xor g115 (n_113, n_222, A[5]);
  nand g116 (n_223, A[3], A[2]);
  nand g117 (n_224, A[5], A[2]);
  nand g118 (n_225, A[3], A[5]);
  nand g119 (n_117, n_223, n_224, n_225);
  xor g120 (n_226, A[0], n_111);
  xor g121 (n_115, n_226, n_112);
  nand g122 (n_227, A[0], n_111);
  nand g123 (n_228, n_112, n_111);
  nand g124 (n_229, A[0], n_112);
  nand g125 (n_120, n_227, n_228, n_229);
  xor g126 (n_230, n_113, n_114);
  xor g127 (n_63, n_230, n_115);
  nand g128 (n_231, n_113, n_114);
  nand g129 (n_232, n_115, n_114);
  nand g130 (n_233, n_113, n_115);
  nand g131 (n_34, n_231, n_232, n_233);
  xor g132 (n_234, A[11], A[8]);
  xor g133 (n_118, n_234, A[4]);
  nand g134 (n_235, A[11], A[8]);
  nand g135 (n_236, A[4], A[8]);
  nand g136 (n_237, A[11], A[4]);
  nand g137 (n_123, n_235, n_236, n_237);
  xor g144 (n_242, n_116, n_117);
  xor g145 (n_121, n_242, n_118);
  nand g146 (n_243, n_116, n_117);
  nand g147 (n_244, n_118, n_117);
  nand g148 (n_245, n_116, n_118);
  nand g149 (n_127, n_243, n_244, n_245);
  xor g150 (n_246, n_67, n_120);
  xor g151 (n_62, n_246, n_121);
  nand g152 (n_247, n_67, n_120);
  nand g153 (n_248, n_121, n_120);
  nand g154 (n_249, n_67, n_121);
  nand g155 (n_33, n_247, n_248, n_249);
  xor g156 (n_250, A[12], A[9]);
  xor g157 (n_124, n_250, A[5]);
  nand g158 (n_251, A[12], A[9]);
  nand g159 (n_252, A[5], A[9]);
  nand g160 (n_253, A[12], A[5]);
  nand g161 (n_42, n_251, n_252, n_253);
  xor g163 (n_125, n_103, A[2]);
  nand g165 (n_256, A[2], A[7]);
  nand g166 (n_257, A[4], A[2]);
  xor g168 (n_258, n_38, n_123);
  xor g169 (n_126, n_258, n_124);
  nand g170 (n_259, n_38, n_123);
  nand g171 (n_260, n_124, n_123);
  nand g172 (n_261, n_38, n_124);
  nand g173 (n_128, n_259, n_260, n_261);
  xor g174 (n_262, n_125, n_126);
  xor g175 (n_61, n_262, n_127);
  nand g176 (n_263, n_125, n_126);
  nand g177 (n_264, n_127, n_126);
  nand g178 (n_265, n_125, n_127);
  nand g179 (n_32, n_263, n_264, n_265);
  xor g180 (n_266, A[13], A[10]);
  xor g181 (n_43, n_266, A[6]);
  nand g182 (n_267, A[13], A[10]);
  nand g183 (n_268, A[6], A[10]);
  nand g184 (n_269, A[13], A[6]);
  nand g185 (n_130, n_267, n_268, n_269);
  xor g187 (n_44, n_104, A[3]);
  nand g189 (n_272, A[3], A[8]);
  xor g192 (n_274, n_41, n_42);
  xor g193 (n_45, n_274, n_43);
  nand g194 (n_275, n_41, n_42);
  nand g195 (n_276, n_43, n_42);
  nand g196 (n_277, n_41, n_43);
  nand g197 (n_134, n_275, n_276, n_277);
  xor g198 (n_278, n_44, n_45);
  xor g199 (n_60, n_278, n_128);
  nand g200 (n_279, n_44, n_45);
  nand g201 (n_280, n_128, n_45);
  nand g202 (n_281, n_44, n_128);
  nand g203 (n_31, n_279, n_280, n_281);
  xor g204 (n_282, A[14], A[11]);
  xor g205 (n_131, n_282, A[7]);
  nand g206 (n_283, A[14], A[11]);
  nand g207 (n_284, A[7], A[11]);
  nand g208 (n_285, A[14], A[7]);
  nand g209 (n_136, n_283, n_284, n_285);
  xor g211 (n_132, n_210, A[4]);
  nand g213 (n_288, A[4], A[9]);
  nand g214 (n_289, A[6], A[4]);
  nand g215 (n_135, n_211, n_288, n_289);
  xor g216 (n_290, n_129, n_130);
  xor g217 (n_133, n_290, n_131);
  nand g218 (n_291, n_129, n_130);
  nand g219 (n_292, n_131, n_130);
  nand g220 (n_293, n_129, n_131);
  nand g221 (n_140, n_291, n_292, n_293);
  xor g222 (n_294, n_132, n_133);
  xor g223 (n_59, n_294, n_134);
  nand g224 (n_295, n_132, n_133);
  nand g225 (n_296, n_134, n_133);
  nand g226 (n_297, n_132, n_134);
  nand g227 (n_30, n_295, n_296, n_297);
  xor g228 (n_298, A[15], A[12]);
  xor g229 (n_137, n_298, A[8]);
  nand g230 (n_299, A[15], A[12]);
  nand g231 (n_300, A[8], A[12]);
  nand g232 (n_301, A[15], A[8]);
  nand g233 (n_143, n_299, n_300, n_301);
  xor g235 (n_138, n_111, A[5]);
  nand g237 (n_304, A[5], A[10]);
  nand g238 (n_305, A[7], A[5]);
  xor g240 (n_306, n_135, n_136);
  xor g241 (n_139, n_306, n_137);
  nand g242 (n_307, n_135, n_136);
  nand g243 (n_308, n_137, n_136);
  nand g244 (n_309, n_135, n_137);
  nand g245 (n_69, n_307, n_308, n_309);
  xor g246 (n_310, n_138, n_139);
  xor g247 (n_58, n_310, n_140);
  nand g248 (n_311, n_138, n_139);
  nand g249 (n_312, n_140, n_139);
  nand g250 (n_313, n_138, n_140);
  nand g251 (n_29, n_311, n_312, n_313);
  xor g254 (n_314, A[9], A[8]);
  xor g255 (n_145, n_314, A[11]);
  nand g256 (n_315, A[9], A[8]);
  nand g258 (n_317, A[9], A[11]);
  nand g259 (n_150, n_315, n_235, n_317);
  nand g264 (n_321, A[6], n_142);
  xor g266 (n_322, n_143, n_144);
  xor g267 (n_147, n_322, n_145);
  nand g268 (n_323, n_143, n_144);
  nand g269 (n_324, n_145, n_144);
  nand g270 (n_325, n_143, n_145);
  nand g271 (n_154, n_323, n_324, n_325);
  xor g272 (n_326, n_146, n_147);
  xor g273 (n_57, n_326, n_69);
  nand g274 (n_327, n_146, n_147);
  nand g275 (n_328, n_69, n_147);
  nand g276 (n_329, n_146, n_69);
  nand g277 (n_28, n_327, n_328, n_329);
  xor g278 (n_148, A[14], A[12]);
  and g279 (n_158, A[14], A[12]);
  xor g280 (n_330, A[9], A[7]);
  xor g281 (n_151, n_330, A[10]);
  nand g282 (n_331, A[9], A[7]);
  nand g284 (n_333, A[9], A[10]);
  nand g289 (n_336, n_149, n_148);
  xor g292 (n_338, n_150, n_151);
  xor g293 (n_155, n_338, n_152);
  nand g294 (n_339, n_150, n_151);
  nand g295 (n_340, n_152, n_151);
  nand g296 (n_341, n_150, n_152);
  nand g297 (n_164, n_339, n_340, n_341);
  xor g298 (n_342, n_153, n_154);
  xor g299 (n_56, n_342, n_155);
  nand g300 (n_343, n_153, n_154);
  nand g301 (n_344, n_155, n_154);
  nand g302 (n_345, n_153, n_155);
  nand g303 (n_27, n_343, n_344, n_345);
  xor g304 (n_157, A[15], A[13]);
  and g305 (n_165, A[15], A[13]);
  xor g306 (n_346, A[10], A[8]);
  xor g307 (n_160, n_346, A[11]);
  nand g308 (n_347, A[10], A[8]);
  nand g310 (n_349, A[10], A[11]);
  nand g311 (n_166, n_347, n_235, n_349);
  nand g315 (n_352, n_158, n_157);
  xor g318 (n_354, n_159, n_160);
  xor g319 (n_163, n_354, n_161);
  nand g320 (n_355, n_159, n_160);
  nand g321 (n_356, n_161, n_160);
  nand g322 (n_357, n_159, n_161);
  nand g323 (n_171, n_355, n_356, n_357);
  xor g324 (n_358, n_162, n_163);
  xor g325 (n_55, n_358, n_164);
  nand g326 (n_359, n_162, n_163);
  nand g327 (n_360, n_164, n_163);
  nand g328 (n_361, n_162, n_164);
  nand g329 (n_26, n_359, n_360, n_361);
  xor g331 (n_167, n_362, A[11]);
  nand g335 (n_174, n_363, n_283, n_365);
  xor g337 (n_169, n_250, n_165);
  nand g339 (n_368, n_165, A[12]);
  nand g340 (n_369, A[9], n_165);
  nand g341 (n_176, n_251, n_368, n_369);
  xor g342 (n_370, n_166, n_167);
  xor g343 (n_170, n_370, n_168);
  nand g344 (n_371, n_166, n_167);
  nand g345 (n_372, n_168, n_167);
  nand g346 (n_373, n_166, n_168);
  nand g347 (n_178, n_371, n_372, n_373);
  xor g348 (n_374, n_169, n_170);
  xor g349 (n_54, n_374, n_171);
  nand g350 (n_375, n_169, n_170);
  nand g351 (n_376, n_171, n_170);
  nand g352 (n_377, n_169, n_171);
  nand g353 (n_25, n_375, n_376, n_377);
  nand g360 (n_381, A[10], A[12]);
  xor g362 (n_382, n_157, n_174);
  xor g363 (n_177, n_382, n_175);
  nand g364 (n_383, n_157, n_174);
  nand g365 (n_384, n_175, n_174);
  nand g366 (n_385, n_157, n_175);
  nand g367 (n_183, n_383, n_384, n_385);
  xor g368 (n_386, n_176, n_177);
  xor g369 (n_53, n_386, n_178);
  nand g370 (n_387, n_176, n_177);
  nand g371 (n_388, n_178, n_177);
  nand g372 (n_389, n_176, n_178);
  nand g373 (n_52, n_387, n_388, n_389);
  xor g380 (n_394, A[13], n_165);
  xor g381 (n_182, n_394, n_180);
  nand g382 (n_395, A[13], n_165);
  nand g383 (n_396, n_180, n_165);
  nand g384 (n_397, A[13], n_180);
  nand g385 (n_188, n_395, n_396, n_397);
  xor g386 (n_398, n_167, n_182);
  xor g387 (n_24, n_398, n_183);
  nand g388 (n_399, n_167, n_182);
  nand g389 (n_400, n_183, n_182);
  nand g390 (n_401, n_167, n_183);
  nand g391 (n_51, n_399, n_400, n_401);
  xor g392 (n_185, A[15], A[14]);
  and g393 (n_189, A[15], A[14]);
  nand g397 (n_404, n_185, A[12]);
  xor g400 (n_406, n_174, n_187);
  xor g401 (n_23, n_406, n_188);
  nand g402 (n_407, n_174, n_187);
  nand g403 (n_408, n_188, n_187);
  nand g404 (n_409, n_174, n_188);
  nand g405 (n_50, n_407, n_408, n_409);
  xor g407 (n_190, n_410, A[13]);
  xor g412 (n_414, n_189, n_190);
  xor g413 (n_22, n_414, n_191);
  nand g414 (n_415, n_189, n_190);
  nand g415 (n_416, n_191, n_190);
  nand g416 (n_417, n_189, n_191);
  nand g417 (n_49, n_415, n_416, n_417);
  xor g419 (n_21, n_362, n_192);
  nand g421 (n_420, n_192, A[14]);
  nand g423 (n_48, n_363, n_420, n_421);
  xor g26 (Z[3], A[3], A[0]);
  nand g31 (n_448, n_215, n_445, n_446);
  nand g34 (n_449, A[2], n_68);
  nand g35 (n_450, A[2], n_448);
  nand g36 (n_451, n_68, n_448);
  nand g37 (n_453, n_449, n_450, n_451);
  xor g38 (n_452, A[2], n_68);
  xor g39 (Z[5], n_448, n_452);
  nand g40 (n_454, n_39, n_67);
  nand g41 (n_455, n_39, n_453);
  nand g42 (n_456, n_67, n_453);
  nand g43 (n_458, n_454, n_455, n_456);
  xor g44 (n_457, n_39, n_67);
  xor g45 (Z[6], n_453, n_457);
  nand g46 (n_459, n_38, n_66);
  nand g47 (n_460, n_38, n_458);
  nand g48 (n_461, n_66, n_458);
  nand g49 (n_463, n_459, n_460, n_461);
  xor g50 (n_462, n_38, n_66);
  xor g51 (Z[7], n_458, n_462);
  nand g52 (n_464, n_37, n_65);
  nand g53 (n_465, n_37, n_463);
  nand g54 (n_466, n_65, n_463);
  nand g55 (n_468, n_464, n_465, n_466);
  xor g56 (n_467, n_37, n_65);
  xor g57 (Z[8], n_463, n_467);
  nand g58 (n_469, n_36, n_64);
  nand g59 (n_470, n_36, n_468);
  nand g60 (n_471, n_64, n_468);
  nand g61 (n_473, n_469, n_470, n_471);
  xor g62 (n_472, n_36, n_64);
  xor g63 (Z[9], n_468, n_472);
  nand g64 (n_474, n_35, n_63);
  nand g65 (n_475, n_35, n_473);
  nand g66 (n_476, n_63, n_473);
  nand g67 (n_478, n_474, n_475, n_476);
  xor g68 (n_477, n_35, n_63);
  xor g431 (Z[10], n_473, n_477);
  nand g432 (n_479, n_34, n_62);
  nand g433 (n_480, n_34, n_478);
  nand g434 (n_481, n_62, n_478);
  nand g435 (n_483, n_479, n_480, n_481);
  xor g436 (n_482, n_34, n_62);
  xor g437 (Z[11], n_478, n_482);
  nand g438 (n_484, n_33, n_61);
  nand g439 (n_485, n_33, n_483);
  nand g440 (n_486, n_61, n_483);
  nand g441 (n_488, n_484, n_485, n_486);
  xor g442 (n_487, n_33, n_61);
  xor g443 (Z[12], n_483, n_487);
  nand g444 (n_489, n_32, n_60);
  nand g445 (n_490, n_32, n_488);
  nand g446 (n_491, n_60, n_488);
  nand g447 (n_493, n_489, n_490, n_491);
  xor g448 (n_492, n_32, n_60);
  xor g449 (Z[13], n_488, n_492);
  nand g450 (n_494, n_31, n_59);
  nand g451 (n_495, n_31, n_493);
  nand g452 (n_496, n_59, n_493);
  nand g453 (n_498, n_494, n_495, n_496);
  xor g454 (n_497, n_31, n_59);
  xor g455 (Z[14], n_493, n_497);
  nand g456 (n_499, n_30, n_58);
  nand g457 (n_500, n_30, n_498);
  nand g458 (n_501, n_58, n_498);
  nand g459 (n_503, n_499, n_500, n_501);
  xor g460 (n_502, n_30, n_58);
  xor g461 (Z[15], n_498, n_502);
  nand g462 (n_504, n_29, n_57);
  nand g463 (n_505, n_29, n_503);
  nand g464 (n_506, n_57, n_503);
  nand g465 (n_508, n_504, n_505, n_506);
  xor g466 (n_507, n_29, n_57);
  xor g467 (Z[16], n_503, n_507);
  nand g468 (n_509, n_28, n_56);
  nand g469 (n_510, n_28, n_508);
  nand g470 (n_511, n_56, n_508);
  nand g471 (n_513, n_509, n_510, n_511);
  xor g472 (n_512, n_28, n_56);
  xor g473 (Z[17], n_508, n_512);
  nand g474 (n_514, n_27, n_55);
  nand g475 (n_515, n_27, n_513);
  nand g476 (n_516, n_55, n_513);
  nand g477 (n_518, n_514, n_515, n_516);
  xor g478 (n_517, n_27, n_55);
  xor g479 (Z[18], n_513, n_517);
  nand g480 (n_519, n_26, n_54);
  nand g481 (n_520, n_26, n_518);
  nand g482 (n_521, n_54, n_518);
  nand g483 (n_523, n_519, n_520, n_521);
  xor g484 (n_522, n_26, n_54);
  xor g485 (Z[19], n_518, n_522);
  nand g486 (n_524, n_25, n_53);
  nand g487 (n_525, n_25, n_523);
  nand g488 (n_526, n_53, n_523);
  nand g489 (n_528, n_524, n_525, n_526);
  xor g490 (n_527, n_25, n_53);
  xor g491 (Z[20], n_523, n_527);
  nand g492 (n_529, n_24, n_52);
  nand g493 (n_530, n_24, n_528);
  nand g494 (n_531, n_52, n_528);
  nand g495 (n_533, n_529, n_530, n_531);
  xor g496 (n_532, n_24, n_52);
  xor g497 (Z[21], n_528, n_532);
  nand g498 (n_534, n_23, n_51);
  nand g499 (n_535, n_23, n_533);
  nand g500 (n_536, n_51, n_533);
  nand g501 (n_538, n_534, n_535, n_536);
  xor g502 (n_537, n_23, n_51);
  xor g503 (Z[22], n_533, n_537);
  nand g504 (n_539, n_22, n_50);
  nand g505 (n_540, n_22, n_538);
  nand g506 (n_541, n_50, n_538);
  nand g507 (n_543, n_539, n_540, n_541);
  xor g508 (n_542, n_22, n_50);
  xor g509 (Z[23], n_538, n_542);
  nand g510 (n_544, n_21, n_49);
  nand g511 (n_545, n_21, n_543);
  nand g512 (n_546, n_49, n_543);
  nand g513 (n_548, n_544, n_545, n_546);
  xor g514 (n_547, n_21, n_49);
  xor g515 (Z[24], n_543, n_547);
  nand g518 (n_551, n_48, n_548);
  nand g519 (n_553, n_549, n_550, n_551);
  xor g521 (Z[25], n_548, n_552);
  nand g524 (n_556, A[15], n_553);
  nand g525 (n_558, n_411, n_555, n_556);
  xor g527 (Z[26], n_553, n_410);
  or g538 (n_41, wc, wc0, n_105);
  not gc0 (wc0, n_256);
  not gc (wc, n_257);
  or g539 (n_129, wc1, wc2, n_107);
  not gc2 (wc2, n_225);
  not gc1 (wc1, n_272);
  or g540 (n_144, wc3, wc4, n_116);
  not gc4 (wc4, n_304);
  not gc3 (wc3, n_305);
  xnor g541 (n_142, A[16], A[13]);
  and g542 (n_149, A[13], wc5);
  not gc5 (wc5, A[16]);
  or g543 (n_159, wc6, wc7, n_116);
  not gc7 (wc7, n_331);
  not gc6 (wc6, n_333);
  xnor g547 (n_362, A[16], A[14]);
  or g548 (n_363, wc8, A[16]);
  not gc8 (wc8, A[14]);
  or g549 (n_365, wc9, A[16]);
  not gc9 (wc9, A[11]);
  xnor g550 (n_175, A[12], A[10]);
  or g551 (n_180, A[10], A[12], wc10);
  not gc10 (wc10, n_381);
  xnor g552 (n_187, n_185, A[12]);
  xnor g554 (n_410, A[16], A[15]);
  or g555 (n_411, wc11, A[16]);
  not gc11 (wc11, A[15]);
  xnor g557 (n_146, n_142, A[6]);
  xnor g559 (n_153, n_148, n_149);
  xnor g560 (n_162, n_158, n_157);
  or g561 (n_168, wc12, n_157, n_158);
  not gc12 (wc12, n_352);
  or g562 (n_191, A[12], wc13, n_185);
  not gc13 (wc13, n_404);
  or g563 (n_192, wc14, n_149, n_165);
  not gc14 (wc14, n_411);
  or g564 (n_152, A[6], n_142, wc15);
  not gc15 (wc15, n_321);
  or g565 (n_161, n_149, wc16, n_148);
  not gc16 (wc16, n_336);
  or g566 (n_421, A[16], wc17);
  not gc17 (wc17, n_192);
  or g567 (n_549, A[15], wc18);
  not gc18 (wc18, n_48);
  xnor g568 (n_552, n_48, A[15]);
  or g570 (n_445, wc19, n_204);
  not gc19 (wc19, A[4]);
  or g571 (n_446, wc20, n_204);
  not gc20 (wc20, A[1]);
  xnor g572 (Z[4], n_204, n_214);
  or g573 (n_550, A[15], wc21);
  not gc21 (wc21, n_548);
  or g574 (n_555, A[16], wc22);
  not gc22 (wc22, n_553);
  not g575 (Z[27], n_558);
endmodule

module mult_signed_const_241_GENERIC(A, Z);
  input [16:0] A;
  output [27:0] Z;
  wire [16:0] A;
  wire [27:0] Z;
  mult_signed_const_241_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_308_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * -10357;"
  input [16:0] A;
  output [31:0] Z;
  wire [16:0] A;
  wire [31:0] Z;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_43, n_44, n_45, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_122, n_124, n_125, n_127, n_128, n_130, n_131;
  wire n_134, n_135, n_136, n_138, n_139, n_140, n_141, n_143;
  wire n_144, n_146, n_147, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_156, n_157, n_158, n_159, n_160, n_161, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_187, n_188, n_190, n_191, n_192;
  wire n_194, n_195, n_196, n_197, n_198, n_200, n_201, n_202;
  wire n_203, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_213, n_214, n_216, n_219, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_273, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_292, n_293, n_294, n_295, n_296;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_308, n_309, n_310, n_311, n_312, n_313, n_315, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_357, n_358, n_361, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_413, n_415, n_416, n_417, n_418, n_421, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_430, n_431, n_432, n_433;
  wire n_434, n_437, n_441, n_445, n_449, n_450, n_459, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567;
  wire n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575;
  wire n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591;
  wire n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599;
  wire n_600, n_601, n_602;
  assign Z[0] = A[0];
  assign Z[30] = Z[31];
  xor g91 (n_77, n_223, A[0]);
  nand g95 (n_44, n_224, n_225, n_226);
  xor g97 (n_76, n_227, A[1]);
  nand g101 (n_43, n_228, n_229, n_230);
  xor g103 (n_75, n_231, A[2]);
  nand g107 (n_122, n_232, n_233, n_234);
  nand g113 (n_124, n_236, A[5], A[7]);
  xor g115 (n_74, n_239, n_122);
  nand g117 (n_241, n_122, A[3]);
  nand g119 (n_41, n_240, n_241, n_242);
  nand g125 (n_127, n_244, n_245, n_246);
  xor g126 (n_247, A[4], n_124);
  xor g127 (n_73, n_247, n_125);
  nand g128 (n_248, A[4], n_124);
  nand g129 (n_249, n_125, n_124);
  nand g130 (n_250, A[4], n_125);
  nand g131 (n_40, n_248, n_249, n_250);
  nand g137 (n_130, n_252, n_253, n_254);
  xor g138 (n_255, A[5], n_127);
  xor g139 (n_72, n_255, n_128);
  nand g140 (n_256, A[5], n_127);
  nand g141 (n_257, n_128, n_127);
  nand g142 (n_258, A[5], n_128);
  nand g143 (n_39, n_256, n_257, n_258);
  nand g149 (n_134, n_260, n_261, n_262);
  xor g150 (n_263, A[6], n_130);
  xor g151 (n_71, n_263, n_131);
  nand g152 (n_264, A[6], n_130);
  nand g153 (n_265, n_131, n_130);
  nand g154 (n_266, A[6], n_131);
  nand g155 (n_38, n_264, n_265, n_266);
  nand g161 (n_139, n_268, n_269, n_270);
  xor g163 (n_135, A[0], A[7]);
  xor g168 (n_275, n_134, n_135);
  xor g169 (n_70, n_275, n_136);
  nand g170 (n_276, n_134, n_135);
  nand g171 (n_277, n_136, n_135);
  nand g172 (n_278, n_134, n_136);
  nand g173 (n_37, n_276, n_277, n_278);
  nand g179 (n_143, n_280, n_281, n_282);
  xor g181 (n_141, n_283, n_138);
  nand g183 (n_285, n_138, A[8]);
  nand g185 (n_146, n_284, n_285, n_286);
  xor g186 (n_287, n_139, n_140);
  xor g187 (n_69, n_287, n_141);
  nand g188 (n_288, n_139, n_140);
  nand g189 (n_289, n_141, n_140);
  nand g190 (n_290, n_139, n_141);
  nand g191 (n_36, n_288, n_289, n_290);
  nand g197 (n_150, n_292, n_293, n_294);
  xor g205 (n_147, n_299, n_144);
  nand g207 (n_301, n_144, n_143);
  nand g209 (n_154, n_300, n_301, n_302);
  xor g211 (n_68, n_303, n_147);
  nand g213 (n_305, n_147, n_146);
  nand g215 (n_35, n_304, n_305, n_306);
  nand g221 (n_157, n_308, n_309, n_310);
  xor g228 (n_315, n_149, n_150);
  xor g229 (n_153, n_315, n_151);
  nand g230 (n_316, n_149, n_150);
  nand g231 (n_317, n_151, n_150);
  nand g232 (n_318, n_149, n_151);
  nand g233 (n_161, n_316, n_317, n_318);
  xor g234 (n_319, n_152, n_153);
  xor g235 (n_67, n_319, n_154);
  nand g236 (n_320, n_152, n_153);
  nand g237 (n_321, n_154, n_153);
  nand g238 (n_322, n_152, n_154);
  nand g239 (n_34, n_320, n_321, n_322);
  nand g245 (n_164, n_324, n_325, n_326);
  nand g251 (n_165, n_328, n_329, n_224);
  xor g252 (n_331, n_156, n_157);
  xor g253 (n_160, n_331, n_158);
  nand g254 (n_332, n_156, n_157);
  nand g255 (n_333, n_158, n_157);
  nand g256 (n_334, n_156, n_158);
  nand g257 (n_169, n_332, n_333, n_334);
  xor g258 (n_335, n_159, n_160);
  xor g259 (n_66, n_335, n_161);
  nand g260 (n_336, n_159, n_160);
  nand g261 (n_337, n_161, n_160);
  nand g262 (n_338, n_159, n_161);
  nand g263 (n_33, n_336, n_337, n_338);
  xor g267 (n_166, n_339, A[12]);
  nand g271 (n_173, n_340, n_341, n_342);
  nand g277 (n_175, A[3], n_345, n_346);
  xor g278 (n_347, n_164, n_165);
  xor g279 (n_168, n_347, n_166);
  nand g280 (n_348, n_164, n_165);
  nand g281 (n_349, n_166, n_165);
  nand g282 (n_350, n_164, n_166);
  nand g283 (n_177, n_348, n_349, n_350);
  xor g284 (n_351, n_167, n_168);
  xor g285 (n_65, n_351, n_169);
  nand g286 (n_352, n_167, n_168);
  nand g287 (n_353, n_169, n_168);
  nand g288 (n_354, n_167, n_169);
  nand g289 (n_32, n_352, n_353, n_354);
  nand g297 (n_180, n_232, n_357, n_358);
  xor g299 (n_176, n_219, n_172);
  xor g304 (n_363, n_173, n_174);
  xor g305 (n_178, n_363, n_175);
  nand g306 (n_364, n_173, n_174);
  nand g307 (n_365, n_175, n_174);
  nand g308 (n_366, n_173, n_175);
  nand g309 (n_185, n_364, n_365, n_366);
  xor g310 (n_367, n_176, n_177);
  xor g311 (n_64, n_367, n_178);
  nand g312 (n_368, n_176, n_177);
  nand g313 (n_369, n_178, n_177);
  nand g314 (n_370, n_176, n_178);
  nand g315 (n_31, n_368, n_369, n_370);
  xor g316 (n_345, A[16], A[14]);
  nand g318 (n_372, A[16], A[14]);
  nand g321 (n_188, n_372, n_373, n_374);
  xor g323 (n_183, n_375, n_179);
  nand g327 (n_190, n_376, n_377, n_378);
  xor g328 (n_379, n_180, n_181);
  xor g329 (n_184, n_379, n_182);
  nand g330 (n_380, n_180, n_181);
  nand g331 (n_381, n_182, n_181);
  nand g332 (n_382, n_180, n_182);
  nand g333 (n_192, n_380, n_381, n_382);
  xor g334 (n_383, n_183, n_184);
  xor g335 (n_63, n_383, n_185);
  nand g336 (n_384, n_183, n_184);
  nand g337 (n_385, n_185, n_184);
  nand g338 (n_386, n_183, n_185);
  nand g339 (n_30, n_384, n_385, n_386);
  nand g347 (n_195, A[6], A[8], n_244);
  xor g348 (n_391, n_187, n_188);
  nand g350 (n_392, n_187, n_188);
  nand g353 (n_198, n_392, n_393, n_394);
  xor g354 (n_395, n_190, n_191);
  xor g355 (n_62, n_395, n_192);
  nand g356 (n_396, n_190, n_191);
  nand g357 (n_397, n_192, n_191);
  nand g358 (n_398, n_190, n_192);
  nand g359 (n_61, n_396, n_397, n_398);
  nand g365 (n_201, n_400, n_401, n_402);
  xor g367 (n_197, n_403, n_195);
  nand g369 (n_405, n_195, n_194);
  nand g371 (n_203, n_404, n_405, n_406);
  xor g372 (n_407, n_196, n_197);
  xor g373 (n_29, n_407, n_198);
  nand g374 (n_408, n_196, n_197);
  nand g375 (n_409, n_198, n_197);
  nand g376 (n_410, n_196, n_198);
  nand g377 (n_60, n_408, n_409, n_410);
  xor g381 (n_202, A[8], n_200);
  xor g386 (n_415, n_201, n_202);
  xor g387 (n_28, n_415, n_203);
  nand g388 (n_416, n_201, n_202);
  nand g389 (n_417, n_203, n_202);
  nand g390 (n_418, n_201, n_203);
  nand g391 (n_27, n_416, n_417, n_418);
  xor g395 (n_207, A[9], n_205);
  xor g400 (n_423, n_206, n_207);
  xor g401 (n_59, n_423, n_208);
  nand g402 (n_424, n_206, n_207);
  nand g403 (n_425, n_208, n_207);
  nand g404 (n_426, n_206, n_208);
  nand g405 (n_26, n_424, n_425, n_426);
  nand g411 (n_214, n_428, n_280, n_430);
  xor g412 (n_431, n_209, n_210);
  xor g413 (n_58, n_431, n_211);
  nand g414 (n_432, n_209, n_210);
  nand g415 (n_433, n_211, n_210);
  nand g416 (n_434, n_209, n_211);
  nand g417 (n_57, n_432, n_433, n_434);
  nand g423 (n_437, n_214, n_213);
  nand g19 (n_467, n_463, n_464, n_465);
  nand g24 (n_470, n_78, n_467);
  nand g25 (n_472, n_468, n_469, n_470);
  xor g27 (Z[3], n_467, n_471);
  nand g28 (n_473, n_45, n_77);
  nand g29 (n_474, n_45, n_472);
  nand g30 (n_475, n_77, n_472);
  nand g31 (n_477, n_473, n_474, n_475);
  xor g32 (n_476, n_45, n_77);
  xor g33 (Z[4], n_472, n_476);
  nand g34 (n_478, n_44, n_76);
  nand g35 (n_479, n_44, n_477);
  nand g36 (n_480, n_76, n_477);
  nand g37 (n_482, n_478, n_479, n_480);
  xor g38 (n_481, n_44, n_76);
  xor g39 (Z[5], n_477, n_481);
  nand g40 (n_483, n_43, n_75);
  nand g41 (n_484, n_43, n_482);
  nand g42 (n_485, n_75, n_482);
  nand g43 (n_487, n_483, n_484, n_485);
  xor g44 (n_486, n_43, n_75);
  xor g45 (Z[6], n_482, n_486);
  nand g48 (n_490, n_74, n_487);
  nand g49 (n_492, n_488, n_489, n_490);
  xor g51 (Z[7], n_487, n_491);
  nand g52 (n_493, n_41, n_73);
  nand g53 (n_494, n_41, n_492);
  nand g54 (n_495, n_73, n_492);
  nand g55 (n_497, n_493, n_494, n_495);
  xor g56 (n_496, n_41, n_73);
  xor g57 (Z[8], n_492, n_496);
  nand g58 (n_498, n_40, n_72);
  nand g59 (n_499, n_40, n_497);
  nand g60 (n_500, n_72, n_497);
  nand g61 (n_502, n_498, n_499, n_500);
  xor g62 (n_501, n_40, n_72);
  xor g63 (Z[9], n_497, n_501);
  nand g64 (n_503, n_39, n_71);
  nand g65 (n_504, n_39, n_502);
  nand g66 (n_505, n_71, n_502);
  nand g67 (n_507, n_503, n_504, n_505);
  xor g68 (n_506, n_39, n_71);
  xor g69 (Z[10], n_502, n_506);
  nand g70 (n_508, n_38, n_70);
  nand g71 (n_509, n_38, n_507);
  nand g72 (n_510, n_70, n_507);
  nand g73 (n_512, n_508, n_509, n_510);
  xor g74 (n_511, n_38, n_70);
  xor g75 (Z[11], n_507, n_511);
  nand g76 (n_513, n_37, n_69);
  nand g77 (n_514, n_37, n_512);
  nand g78 (n_515, n_69, n_512);
  nand g79 (n_517, n_513, n_514, n_515);
  xor g80 (n_516, n_37, n_69);
  xor g81 (Z[12], n_512, n_516);
  nand g82 (n_518, n_36, n_68);
  nand g83 (n_519, n_36, n_517);
  nand g84 (n_520, n_68, n_517);
  nand g85 (n_522, n_518, n_519, n_520);
  xor g466 (n_521, n_36, n_68);
  xor g467 (Z[13], n_517, n_521);
  nand g468 (n_523, n_35, n_67);
  nand g469 (n_524, n_35, n_522);
  nand g470 (n_525, n_67, n_522);
  nand g471 (n_527, n_523, n_524, n_525);
  xor g472 (n_526, n_35, n_67);
  xor g473 (Z[14], n_522, n_526);
  nand g474 (n_528, n_34, n_66);
  nand g475 (n_529, n_34, n_527);
  nand g476 (n_530, n_66, n_527);
  nand g477 (n_532, n_528, n_529, n_530);
  xor g478 (n_531, n_34, n_66);
  xor g479 (Z[15], n_527, n_531);
  nand g480 (n_533, n_33, n_65);
  nand g481 (n_534, n_33, n_532);
  nand g482 (n_535, n_65, n_532);
  nand g483 (n_537, n_533, n_534, n_535);
  xor g484 (n_536, n_33, n_65);
  xor g485 (Z[16], n_532, n_536);
  nand g486 (n_538, n_32, n_64);
  nand g487 (n_539, n_32, n_537);
  nand g488 (n_540, n_64, n_537);
  nand g489 (n_542, n_538, n_539, n_540);
  xor g490 (n_541, n_32, n_64);
  xor g491 (Z[17], n_537, n_541);
  nand g492 (n_543, n_31, n_63);
  nand g493 (n_544, n_31, n_542);
  nand g494 (n_545, n_63, n_542);
  nand g495 (n_547, n_543, n_544, n_545);
  xor g496 (n_546, n_31, n_63);
  xor g497 (Z[18], n_542, n_546);
  nand g498 (n_548, n_30, n_62);
  nand g499 (n_549, n_30, n_547);
  nand g500 (n_550, n_62, n_547);
  nand g501 (n_552, n_548, n_549, n_550);
  xor g502 (n_551, n_30, n_62);
  xor g503 (Z[19], n_547, n_551);
  nand g504 (n_553, n_29, n_61);
  nand g505 (n_554, n_29, n_552);
  nand g506 (n_555, n_61, n_552);
  nand g507 (n_557, n_553, n_554, n_555);
  xor g508 (n_556, n_29, n_61);
  xor g509 (Z[20], n_552, n_556);
  nand g510 (n_558, n_28, n_60);
  nand g511 (n_559, n_28, n_557);
  nand g512 (n_560, n_60, n_557);
  nand g513 (n_562, n_558, n_559, n_560);
  xor g514 (n_561, n_28, n_60);
  xor g515 (Z[21], n_557, n_561);
  nand g516 (n_563, n_27, n_59);
  nand g517 (n_564, n_27, n_562);
  nand g518 (n_565, n_59, n_562);
  nand g519 (n_567, n_563, n_564, n_565);
  xor g520 (n_566, n_27, n_59);
  xor g521 (Z[22], n_562, n_566);
  nand g522 (n_568, n_26, n_58);
  nand g523 (n_569, n_26, n_567);
  nand g524 (n_570, n_58, n_567);
  nand g525 (n_572, n_568, n_569, n_570);
  xor g526 (n_571, n_26, n_58);
  xor g527 (Z[23], n_567, n_571);
  nand g528 (n_573, n_25, n_57);
  nand g529 (n_574, n_25, n_572);
  nand g530 (n_575, n_57, n_572);
  nand g531 (n_577, n_573, n_574, n_575);
  xor g532 (n_576, n_25, n_57);
  xor g533 (Z[24], n_572, n_576);
  nand g534 (n_578, n_24, n_56);
  nand g535 (n_579, n_24, n_577);
  nand g536 (n_580, n_56, n_577);
  nand g537 (n_582, n_578, n_579, n_580);
  xor g538 (n_581, n_24, n_56);
  xor g539 (Z[25], n_577, n_581);
  nand g540 (n_583, n_23, n_55);
  nand g541 (n_584, n_23, n_582);
  nand g542 (n_585, n_55, n_582);
  nand g543 (n_587, n_583, n_584, n_585);
  xor g544 (n_586, n_23, n_55);
  xor g545 (Z[26], n_582, n_586);
  nand g546 (n_588, n_22, n_54);
  nand g547 (n_589, n_22, n_587);
  nand g548 (n_590, n_54, n_587);
  nand g549 (n_592, n_588, n_589, n_590);
  xor g550 (n_591, n_22, n_54);
  xor g551 (Z[27], n_587, n_591);
  nand g552 (n_593, A[15], n_53);
  nand g553 (n_594, A[15], n_592);
  nand g554 (n_595, n_53, n_592);
  nand g555 (n_597, n_593, n_594, n_595);
  xor g556 (n_596, A[15], n_53);
  xor g557 (Z[28], n_592, n_596);
  nand g559 (n_599, A[16], n_597);
  nand g561 (n_602, n_598, n_599, n_600);
  xor g563 (Z[29], n_597, n_601);
  xor g572 (n_78, A[3], A[1]);
  nor g573 (n_45, A[3], A[1]);
  xor g574 (n_223, A[4], A[2]);
  or g575 (n_224, A[4], A[2]);
  or g576 (n_225, wc, A[2]);
  not gc (wc, A[0]);
  or g577 (n_226, wc0, A[4]);
  not gc0 (wc0, A[0]);
  xor g578 (n_227, A[5], A[3]);
  or g579 (n_228, A[5], A[3]);
  or g580 (n_229, wc1, A[3]);
  not gc1 (wc1, A[1]);
  or g581 (n_230, wc2, A[5]);
  not gc2 (wc2, A[1]);
  xor g582 (n_231, A[6], A[4]);
  or g583 (n_232, A[6], A[4]);
  or g584 (n_233, wc3, A[4]);
  not gc3 (wc3, A[2]);
  or g585 (n_234, wc4, A[6]);
  not gc4 (wc4, A[2]);
  xor g586 (n_235, A[7], A[5]);
  or g587 (n_236, A[7], A[5]);
  xnor g588 (n_239, A[3], A[0]);
  or g589 (n_240, A[0], wc5);
  not gc5 (wc5, A[3]);
  xor g590 (n_243, A[8], A[6]);
  or g591 (n_244, A[8], A[6]);
  or g592 (n_245, A[6], A[1]);
  or g593 (n_246, A[8], A[1]);
  xor g594 (n_251, A[9], A[7]);
  or g595 (n_252, A[9], A[7]);
  or g596 (n_253, A[7], A[2]);
  or g597 (n_254, A[9], A[2]);
  xor g598 (n_259, A[10], A[8]);
  or g599 (n_260, A[10], A[8]);
  or g600 (n_261, A[8], A[3]);
  or g601 (n_262, A[10], A[3]);
  xor g602 (n_267, A[11], A[9]);
  or g603 (n_268, A[11], A[9]);
  or g604 (n_269, A[9], A[4]);
  or g605 (n_270, A[11], A[4]);
  or g606 (n_273, A[0], wc6);
  not gc6 (wc6, A[7]);
  xor g607 (n_279, A[12], A[10]);
  or g608 (n_280, A[12], A[10]);
  or g609 (n_281, A[10], A[5]);
  or g610 (n_282, A[12], A[5]);
  xnor g611 (n_283, A[8], A[1]);
  or g612 (n_284, A[1], wc7);
  not gc7 (wc7, A[8]);
  xor g613 (n_213, A[13], A[11]);
  or g614 (n_292, A[13], A[11]);
  or g615 (n_293, A[11], A[6]);
  or g616 (n_294, A[13], A[6]);
  xnor g617 (n_295, A[9], A[2]);
  or g618 (n_296, A[2], wc8);
  not gc8 (wc8, A[9]);
  xor g619 (n_216, A[14], A[12]);
  or g620 (n_308, A[14], A[12]);
  or g621 (n_309, A[12], A[7]);
  or g622 (n_310, A[14], A[7]);
  xnor g623 (n_311, A[10], A[3]);
  or g624 (n_312, A[3], wc9);
  not gc9 (wc9, A[10]);
  or g625 (n_313, A[1], wc10);
  not gc10 (wc10, A[10]);
  xor g627 (n_219, A[15], A[13]);
  or g628 (n_324, A[15], A[13]);
  or g629 (n_325, A[13], A[8]);
  or g630 (n_326, A[15], A[8]);
  xnor g631 (n_327, A[11], A[4]);
  or g632 (n_328, A[4], wc11);
  not gc11 (wc11, A[11]);
  or g633 (n_329, A[2], wc12);
  not gc12 (wc12, A[11]);
  and g635 (n_172, wc13, A[16]);
  not gc13 (wc13, A[14]);
  xor g636 (n_339, A[9], A[5]);
  or g637 (n_340, A[9], A[5]);
  or g638 (n_341, A[5], wc14);
  not gc14 (wc14, A[12]);
  or g639 (n_342, A[9], wc15);
  not gc15 (wc15, A[12]);
  and g641 (n_179, A[13], wc16);
  not gc16 (wc16, A[15]);
  or g642 (n_357, A[10], A[4]);
  or g643 (n_358, A[10], A[6]);
  xnor g644 (n_181, n_345, A[7]);
  or g645 (n_373, A[7], wc17);
  not gc17 (wc17, A[14]);
  or g646 (n_374, A[7], wc18);
  not gc18 (wc18, A[16]);
  xor g647 (n_375, A[11], A[5]);
  or g648 (n_376, A[11], A[5]);
  xnor g649 (n_187, A[15], A[12]);
  and g650 (n_194, wc19, A[15]);
  not gc19 (wc19, A[12]);
  xor g651 (n_399, A[16], A[13]);
  or g652 (n_400, A[16], A[13]);
  or g653 (n_401, A[13], A[7]);
  or g654 (n_402, A[16], A[7]);
  xor g655 (n_200, A[14], A[10]);
  nor g656 (n_205, A[14], A[10]);
  xor g657 (n_206, A[15], A[11]);
  nor g658 (n_209, A[15], A[11]);
  xnor g659 (n_427, A[16], A[12]);
  or g660 (n_428, A[12], wc20);
  not gc20 (wc20, A[16]);
  or g661 (n_430, A[10], wc21);
  not gc21 (wc21, A[16]);
  xnor g667 (n_125, n_243, A[1]);
  xnor g668 (n_128, n_251, A[2]);
  xnor g669 (n_131, n_259, A[3]);
  xnor g670 (n_136, n_267, A[4]);
  or g671 (n_138, wc22, A[7], wc23);
  not gc23 (wc23, n_273);
  not gc22 (wc22, A[0]);
  xnor g672 (n_140, n_279, A[5]);
  xnor g673 (n_144, n_213, A[6]);
  or g675 (n_149, wc24, A[9], wc25);
  not gc25 (wc25, n_296);
  not gc24 (wc24, A[2]);
  xnor g676 (n_151, n_216, A[7]);
  xnor g677 (n_152, n_311, A[1]);
  or g678 (n_156, wc26, wc27, n_45);
  not gc27 (wc27, n_312);
  not gc26 (wc26, n_313);
  xnor g679 (n_158, n_219, A[8]);
  xnor g680 (n_159, n_327, A[2]);
  xnor g681 (n_167, n_345, A[3]);
  or g682 (n_346, n_345, A[3]);
  xnor g683 (n_174, n_231, A[10]);
  or g684 (n_361, wc28, n_219);
  not gc28 (wc28, n_172);
  or g685 (n_377, A[11], wc29);
  not gc29 (wc29, n_179);
  or g686 (n_378, A[5], wc30);
  not gc30 (wc30, n_179);
  xnor g688 (n_196, n_399, A[7]);
  xnor g689 (n_403, n_194, A[9]);
  or g690 (n_404, A[9], wc31);
  not gc31 (wc31, n_194);
  or g691 (n_413, A[8], wc32);
  not gc32 (wc32, n_200);
  or g693 (n_421, A[9], wc33);
  not gc33 (wc33, n_205);
  xnor g695 (n_210, n_427, A[10]);
  or g698 (n_441, wc34, n_292);
  not gc34 (wc34, n_216);
  or g700 (n_445, wc35, n_308);
  not gc35 (wc35, n_219);
  xor g701 (n_54, n_345, n_324);
  or g702 (n_449, n_324, A[14]);
  or g703 (n_450, wc36, n_324);
  not gc36 (wc36, A[16]);
  or g704 (n_463, A[0], wc37);
  not gc37 (wc37, A[2]);
  xnor g705 (n_466, A[2], A[0]);
  or g706 (n_468, A[2], wc38);
  not gc38 (wc38, n_78);
  xnor g707 (n_471, n_78, A[2]);
  or g708 (n_598, A[15], wc39);
  not gc39 (wc39, A[16]);
  xnor g709 (n_601, A[16], A[15]);
  or g710 (n_242, A[0], wc40);
  not gc40 (wc40, n_122);
  or g711 (n_286, A[1], wc41);
  not gc41 (wc41, n_138);
  xnor g712 (n_299, n_143, A[0]);
  or g713 (n_300, A[0], wc42);
  not gc42 (wc42, n_143);
  or g714 (n_302, A[0], wc43);
  not gc43 (wc43, n_144);
  or g715 (n_182, wc44, n_172, wc45);
  not gc45 (wc45, n_219);
  not gc44 (wc44, n_361);
  or g716 (n_393, n_243, wc46);
  not gc46 (wc46, n_188);
  or g717 (n_394, wc47, n_243);
  not gc47 (wc47, n_187);
  or g718 (n_406, A[9], wc48);
  not gc48 (wc48, n_195);
  or g719 (n_208, wc49, wc50, n_200);
  not gc50 (wc50, n_413);
  not gc49 (wc49, A[8]);
  or g720 (n_211, wc51, wc52, n_205);
  not gc52 (wc52, n_421);
  not gc51 (wc51, A[9]);
  xnor g721 (n_25, n_214, n_213);
  xor g723 (n_56, n_292, n_216);
  or g724 (n_23, wc53, n_216, wc54);
  not gc54 (wc54, n_292);
  not gc53 (wc53, n_441);
  xor g725 (n_55, n_308, n_219);
  or g726 (n_22, wc55, n_219, wc56);
  not gc56 (wc56, n_308);
  not gc55 (wc55, n_445);
  or g727 (n_53, wc57, wc58, n_172);
  not gc58 (wc58, n_449);
  not gc57 (wc57, n_450);
  or g728 (n_459, A[1], A[0]);
  xor g729 (Z[1], A[1], A[0]);
  xnor g730 (n_191, n_391, n_243);
  or g731 (n_24, n_213, wc59, n_214);
  not gc59 (wc59, n_437);
  or g733 (n_488, n_235, wc60);
  not gc60 (wc60, n_74);
  xnor g734 (n_491, n_74, n_235);
  xnor g735 (n_303, n_146, n_295);
  or g736 (n_304, n_295, wc61);
  not gc61 (wc61, n_146);
  or g737 (n_306, n_295, wc62);
  not gc62 (wc62, n_147);
  or g738 (n_464, n_459, A[0]);
  or g739 (n_465, wc63, n_459);
  not gc63 (wc63, A[2]);
  xnor g740 (Z[2], n_466, n_459);
  or g741 (n_469, A[2], wc64);
  not gc64 (wc64, n_467);
  or g742 (n_489, n_235, wc65);
  not gc65 (wc65, n_487);
  or g743 (n_600, A[15], wc66);
  not gc66 (wc66, n_597);
  not g744 (Z[31], n_602);
endmodule

module mult_signed_const_308_GENERIC(A, Z);
  input [16:0] A;
  output [31:0] Z;
  wire [16:0] A;
  wire [31:0] Z;
  mult_signed_const_308_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_403_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 104741;"
  input [16:0] A;
  output [33:0] Z;
  wire [16:0] A;
  wire [33:0] Z;
  wire n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27;
  wire n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_53, n_54;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_83, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_152, n_153, n_154, n_155, n_156, n_157, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_209, n_210, n_212;
  wire n_213, n_214, n_215, n_220, n_221, n_222, n_223, n_224;
  wire n_226, n_228, n_229, n_230, n_231, n_233, n_235, n_236;
  wire n_237, n_238, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_256, n_261, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_343, n_344, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_365, n_366, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_382, n_384, n_387, n_389;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_409, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_427, n_428, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_448, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_467;
  wire n_468, n_469, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_491, n_493, n_494, n_495, n_496, n_497, n_498, n_499;
  wire n_500, n_501, n_503, n_504, n_507, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531;
  wire n_532, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_579, n_587, n_588;
  wire n_601, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g98 (n_80, A[5], A[0]);
  and g2 (n_45, A[5], A[0]);
  xor g99 (n_261, A[6], A[4]);
  xor g100 (n_79, n_261, A[1]);
  nand g3 (n_262, A[6], A[4]);
  nand g101 (n_263, A[1], A[4]);
  nand g102 (n_264, A[6], A[1]);
  nand g103 (n_44, n_262, n_263, n_264);
  xor g104 (n_265, A[7], A[5]);
  xor g105 (n_78, n_265, A[2]);
  nand g106 (n_266, A[7], A[5]);
  nand g4 (n_267, A[2], A[5]);
  nand g107 (n_268, A[7], A[2]);
  nand g108 (n_43, n_266, n_267, n_268);
  xor g109 (n_121, A[8], A[6]);
  and g110 (n_122, A[8], A[6]);
  xor g111 (n_269, A[0], A[3]);
  xor g112 (n_77, n_269, n_121);
  nand g113 (n_270, A[0], A[3]);
  nand g114 (n_271, n_121, A[3]);
  nand g5 (n_272, A[0], n_121);
  nand g6 (n_42, n_270, n_271, n_272);
  xor g115 (n_273, A[9], A[7]);
  xor g116 (n_123, n_273, A[1]);
  nand g117 (n_274, A[9], A[7]);
  nand g118 (n_275, A[1], A[7]);
  nand g119 (n_276, A[9], A[1]);
  nand g120 (n_124, n_274, n_275, n_276);
  xor g121 (n_277, A[4], n_122);
  xor g122 (n_76, n_277, n_123);
  nand g123 (n_278, A[4], n_122);
  nand g124 (n_279, n_123, n_122);
  nand g125 (n_280, A[4], n_123);
  nand g126 (n_41, n_278, n_279, n_280);
  xor g127 (n_281, A[10], A[8]);
  xor g128 (n_125, n_281, A[2]);
  nand g129 (n_282, A[10], A[8]);
  nand g130 (n_283, A[2], A[8]);
  nand g131 (n_284, A[10], A[2]);
  nand g132 (n_127, n_282, n_283, n_284);
  xor g133 (n_285, A[5], n_124);
  xor g134 (n_75, n_285, n_125);
  nand g135 (n_286, A[5], n_124);
  nand g136 (n_287, n_125, n_124);
  nand g137 (n_288, A[5], n_125);
  nand g138 (n_40, n_286, n_287, n_288);
  xor g139 (n_126, A[11], A[9]);
  and g140 (n_130, A[11], A[9]);
  xor g142 (n_128, n_269, A[6]);
  nand g144 (n_291, A[6], A[0]);
  nand g145 (n_292, A[3], A[6]);
  nand g146 (n_131, n_270, n_291, n_292);
  xor g147 (n_293, n_126, n_127);
  xor g148 (n_74, n_293, n_128);
  nand g149 (n_294, n_126, n_127);
  nand g150 (n_295, n_128, n_127);
  nand g151 (n_296, n_126, n_128);
  nand g152 (n_39, n_294, n_295, n_296);
  xor g153 (n_129, A[12], A[10]);
  and g154 (n_134, A[12], A[10]);
  xor g155 (n_297, A[4], A[1]);
  xor g156 (n_132, n_297, A[7]);
  nand g159 (n_300, A[4], A[7]);
  nand g160 (n_135, n_263, n_275, n_300);
  xor g161 (n_301, A[0], n_129);
  xor g162 (n_133, n_301, n_130);
  nand g163 (n_302, A[0], n_129);
  nand g164 (n_303, n_130, n_129);
  nand g165 (n_304, A[0], n_130);
  nand g166 (n_138, n_302, n_303, n_304);
  xor g167 (n_305, n_131, n_132);
  xor g168 (n_73, n_305, n_133);
  nand g169 (n_306, n_131, n_132);
  nand g170 (n_307, n_133, n_132);
  nand g171 (n_308, n_131, n_133);
  nand g172 (n_38, n_306, n_307, n_308);
  xor g173 (n_309, A[13], A[11]);
  xor g174 (n_136, n_309, A[5]);
  nand g175 (n_310, A[13], A[11]);
  nand g176 (n_311, A[5], A[11]);
  nand g177 (n_312, A[13], A[5]);
  nand g178 (n_141, n_310, n_311, n_312);
  xor g179 (n_313, A[2], A[8]);
  xor g180 (n_137, n_313, A[1]);
  nand g182 (n_315, A[1], A[8]);
  nand g183 (n_316, A[2], A[1]);
  nand g184 (n_140, n_283, n_315, n_316);
  xor g185 (n_317, n_134, n_135);
  xor g186 (n_139, n_317, n_136);
  nand g187 (n_318, n_134, n_135);
  nand g188 (n_319, n_136, n_135);
  nand g189 (n_320, n_134, n_136);
  nand g190 (n_145, n_318, n_319, n_320);
  xor g191 (n_321, n_137, n_138);
  xor g192 (n_72, n_321, n_139);
  nand g193 (n_322, n_137, n_138);
  nand g194 (n_323, n_139, n_138);
  nand g195 (n_324, n_137, n_139);
  nand g196 (n_37, n_322, n_323, n_324);
  xor g197 (n_325, A[14], A[12]);
  xor g198 (n_142, n_325, A[6]);
  nand g199 (n_326, A[14], A[12]);
  nand g200 (n_327, A[6], A[12]);
  nand g201 (n_328, A[14], A[6]);
  nand g202 (n_147, n_326, n_327, n_328);
  xor g203 (n_329, A[3], A[9]);
  xor g204 (n_143, n_329, A[2]);
  nand g205 (n_330, A[3], A[9]);
  nand g206 (n_331, A[2], A[9]);
  nand g207 (n_332, A[3], A[2]);
  nand g208 (n_148, n_330, n_331, n_332);
  xor g209 (n_333, n_140, n_141);
  xor g210 (n_144, n_333, n_142);
  nand g211 (n_334, n_140, n_141);
  nand g212 (n_335, n_142, n_141);
  nand g213 (n_336, n_140, n_142);
  nand g214 (n_49, n_334, n_335, n_336);
  xor g215 (n_337, n_143, n_144);
  xor g216 (n_71, n_337, n_145);
  nand g217 (n_338, n_143, n_144);
  nand g218 (n_339, n_145, n_144);
  nand g219 (n_340, n_143, n_145);
  nand g220 (n_36, n_338, n_339, n_340);
  xor g221 (n_146, A[15], A[13]);
  and g222 (n_149, A[15], A[13]);
  xor g223 (n_341, A[7], A[4]);
  xor g224 (n_46, n_341, A[10]);
  nand g226 (n_343, A[10], A[4]);
  nand g227 (n_344, A[7], A[10]);
  nand g228 (n_150, n_300, n_343, n_344);
  xor g230 (n_47, n_269, n_146);
  nand g232 (n_347, n_146, A[0]);
  nand g233 (n_348, A[3], n_146);
  nand g234 (n_154, n_270, n_347, n_348);
  xor g235 (n_349, n_147, n_148);
  xor g236 (n_48, n_349, n_46);
  nand g237 (n_350, n_147, n_148);
  nand g238 (n_351, n_46, n_148);
  nand g239 (n_352, n_147, n_46);
  nand g240 (n_155, n_350, n_351, n_352);
  xor g241 (n_353, n_47, n_48);
  xor g242 (n_70, n_353, n_49);
  nand g243 (n_354, n_47, n_48);
  nand g244 (n_355, n_49, n_48);
  nand g245 (n_356, n_47, n_49);
  nand g246 (n_35, n_354, n_355, n_356);
  xor g248 (n_153, n_357, A[8]);
  nand g250 (n_359, A[8], A[14]);
  nand g252 (n_159, n_358, n_359, n_360);
  xor g259 (n_365, A[11], A[4]);
  xor g260 (n_152, n_365, A[1]);
  nand g261 (n_366, A[11], A[4]);
  nand g263 (n_368, A[11], A[1]);
  nand g264 (n_161, n_366, n_263, n_368);
  xor g265 (n_369, n_149, n_150);
  nand g267 (n_370, n_149, n_150);
  nand g270 (n_165, n_370, n_371, n_372);
  xor g271 (n_373, n_152, n_153);
  xor g272 (n_157, n_373, n_154);
  nand g273 (n_374, n_152, n_153);
  nand g274 (n_375, n_154, n_153);
  nand g275 (n_376, n_152, n_154);
  nand g276 (n_167, n_374, n_375, n_376);
  xor g277 (n_377, n_155, n_156);
  xor g278 (n_69, n_377, n_157);
  nand g279 (n_378, n_155, n_156);
  nand g280 (n_379, n_157, n_156);
  nand g281 (n_380, n_155, n_157);
  nand g282 (n_34, n_378, n_379, n_380);
  xor g283 (n_188, A[15], A[12]);
  xor g284 (n_162, n_188, A[6]);
  nand g285 (n_382, A[15], A[12]);
  nand g287 (n_384, A[15], A[6]);
  nand g288 (n_171, n_382, n_327, n_384);
  nand g292 (n_387, A[9], A[5]);
  xor g295 (n_389, A[2], A[1]);
  xor g296 (n_164, n_389, n_159);
  nand g298 (n_391, n_159, A[1]);
  nand g299 (n_392, A[2], n_159);
  nand g300 (n_174, n_316, n_391, n_392);
  xor g301 (n_393, n_160, n_161);
  xor g302 (n_166, n_393, n_162);
  nand g303 (n_394, n_160, n_161);
  nand g304 (n_395, n_162, n_161);
  nand g305 (n_396, n_160, n_162);
  nand g306 (n_175, n_394, n_395, n_396);
  xor g307 (n_397, n_163, n_164);
  xor g308 (n_168, n_397, n_165);
  nand g309 (n_398, n_163, n_164);
  nand g310 (n_399, n_165, n_164);
  nand g311 (n_400, n_163, n_165);
  nand g312 (n_81, n_398, n_399, n_400);
  xor g313 (n_401, n_166, n_167);
  xor g314 (n_68, n_401, n_168);
  nand g315 (n_402, n_166, n_167);
  nand g316 (n_403, n_168, n_167);
  nand g317 (n_404, n_166, n_168);
  nand g318 (n_33, n_402, n_403, n_404);
  xor g321 (n_405, A[7], A[6]);
  xor g322 (n_172, n_405, A[10]);
  nand g323 (n_406, A[7], A[6]);
  nand g324 (n_407, A[10], A[6]);
  nand g326 (n_179, n_406, n_407, n_344);
  xor g327 (n_409, A[3], A[2]);
  xor g328 (n_173, n_409, n_169);
  nand g330 (n_411, n_169, A[2]);
  nand g331 (n_412, A[3], n_169);
  nand g332 (n_182, n_332, n_411, n_412);
  xor g333 (n_413, n_170, n_171);
  xor g334 (n_176, n_413, n_172);
  nand g335 (n_414, n_170, n_171);
  nand g336 (n_415, n_172, n_171);
  nand g337 (n_416, n_170, n_172);
  nand g338 (n_183, n_414, n_415, n_416);
  xor g339 (n_417, n_173, n_174);
  xor g340 (n_177, n_417, n_175);
  nand g341 (n_418, n_173, n_174);
  nand g342 (n_419, n_175, n_174);
  nand g343 (n_420, n_173, n_175);
  nand g344 (n_186, n_418, n_419, n_420);
  xor g345 (n_421, n_176, n_177);
  xor g346 (n_67, n_421, n_81);
  nand g347 (n_422, n_176, n_177);
  nand g348 (n_423, n_81, n_177);
  nand g349 (n_424, n_176, n_81);
  nand g350 (n_32, n_422, n_423, n_424);
  xor g351 (n_83, A[14], A[11]);
  and g352 (n_189, A[14], A[11]);
  xor g354 (n_180, n_341, A[8]);
  nand g356 (n_427, A[8], A[4]);
  nand g357 (n_428, A[7], A[8]);
  nand g358 (n_190, n_300, n_427, n_428);
  nand g363 (n_432, A[3], n_83);
  xor g365 (n_433, n_178, n_179);
  xor g366 (n_184, n_433, n_180);
  nand g367 (n_434, n_178, n_179);
  nand g368 (n_435, n_180, n_179);
  nand g369 (n_436, n_178, n_180);
  nand g370 (n_194, n_434, n_435, n_436);
  xor g371 (n_437, n_181, n_182);
  xor g372 (n_185, n_437, n_183);
  nand g373 (n_438, n_181, n_182);
  nand g374 (n_439, n_183, n_182);
  nand g375 (n_440, n_181, n_183);
  nand g376 (n_197, n_438, n_439, n_440);
  xor g377 (n_441, n_184, n_185);
  xor g378 (n_66, n_441, n_186);
  nand g379 (n_442, n_184, n_185);
  nand g380 (n_443, n_186, n_185);
  nand g381 (n_444, n_184, n_186);
  nand g382 (n_31, n_442, n_443, n_444);
  xor g385 (n_445, A[8], A[5]);
  xor g386 (n_191, n_445, A[9]);
  nand g387 (n_446, A[8], A[5]);
  nand g389 (n_448, A[8], A[9]);
  nand g390 (n_199, n_446, n_387, n_448);
  nand g395 (n_452, A[4], n_188);
  xor g397 (n_453, n_189, n_190);
  xor g398 (n_195, n_453, n_191);
  nand g399 (n_454, n_189, n_190);
  nand g400 (n_455, n_191, n_190);
  nand g401 (n_456, n_189, n_191);
  nand g402 (n_204, n_454, n_455, n_456);
  xor g403 (n_457, n_192, n_193);
  xor g404 (n_196, n_457, n_194);
  nand g405 (n_458, n_192, n_193);
  nand g406 (n_459, n_194, n_193);
  nand g407 (n_460, n_192, n_194);
  nand g408 (n_206, n_458, n_459, n_460);
  xor g409 (n_461, n_195, n_196);
  xor g410 (n_65, n_461, n_197);
  nand g411 (n_462, n_195, n_196);
  nand g412 (n_463, n_197, n_196);
  nand g413 (n_464, n_195, n_197);
  nand g414 (n_30, n_462, n_463, n_464);
  xor g416 (n_201, n_169, A[9]);
  nand g418 (n_467, A[9], A[13]);
  xor g421 (n_469, A[6], A[10]);
  xor g422 (n_200, n_469, A[5]);
  nand g424 (n_471, A[5], A[10]);
  nand g425 (n_472, A[6], A[5]);
  nand g426 (n_209, n_407, n_471, n_472);
  xor g428 (n_203, n_473, n_200);
  nand g430 (n_475, n_200, n_199);
  nand g432 (n_213, n_474, n_475, n_476);
  xor g433 (n_477, n_201, n_202);
  xor g434 (n_205, n_477, n_203);
  nand g435 (n_478, n_201, n_202);
  nand g436 (n_479, n_203, n_202);
  nand g437 (n_480, n_201, n_203);
  nand g438 (n_215, n_478, n_479, n_480);
  xor g439 (n_481, n_204, n_205);
  xor g440 (n_64, n_481, n_206);
  nand g441 (n_482, n_204, n_205);
  nand g442 (n_483, n_206, n_205);
  nand g443 (n_484, n_204, n_206);
  nand g444 (n_29, n_482, n_483, n_484);
  nand g456 (n_491, n_209, n_83);
  xor g459 (n_493, n_210, n_172);
  xor g460 (n_214, n_493, n_212);
  nand g461 (n_494, n_210, n_172);
  nand g462 (n_495, n_212, n_172);
  nand g463 (n_496, n_210, n_212);
  nand g464 (n_224, n_494, n_495, n_496);
  xor g465 (n_497, n_213, n_214);
  xor g466 (n_63, n_497, n_215);
  nand g467 (n_498, n_213, n_214);
  nand g468 (n_499, n_215, n_214);
  nand g469 (n_500, n_213, n_215);
  nand g470 (n_28, n_498, n_499, n_500);
  xor g473 (n_501, A[8], A[7]);
  xor g474 (n_220, n_501, A[11]);
  nand g476 (n_503, A[11], A[7]);
  nand g477 (n_504, A[8], A[11]);
  nand g478 (n_226, n_428, n_503, n_504);
  nand g482 (n_507, n_189, n_188);
  xor g485 (n_509, n_179, n_220);
  xor g486 (n_223, n_509, n_221);
  nand g487 (n_510, n_179, n_220);
  nand g488 (n_511, n_221, n_220);
  nand g489 (n_512, n_179, n_221);
  nand g490 (n_231, n_510, n_511, n_512);
  xor g491 (n_513, n_222, n_223);
  xor g492 (n_62, n_513, n_224);
  nand g493 (n_514, n_222, n_223);
  nand g494 (n_515, n_224, n_223);
  nand g495 (n_516, n_222, n_224);
  nand g496 (n_27, n_514, n_515, n_516);
  xor g503 (n_521, A[8], A[12]);
  nand g505 (n_522, A[8], A[12]);
  nand g508 (n_236, n_522, n_523, n_524);
  xor g509 (n_525, n_226, n_201);
  xor g510 (n_230, n_525, n_228);
  nand g511 (n_526, n_226, n_201);
  nand g512 (n_527, n_228, n_201);
  nand g513 (n_528, n_226, n_228);
  nand g514 (n_238, n_526, n_527, n_528);
  xor g515 (n_529, n_229, n_230);
  xor g516 (n_61, n_529, n_231);
  nand g517 (n_530, n_229, n_230);
  nand g518 (n_531, n_231, n_230);
  nand g519 (n_532, n_229, n_231);
  nand g520 (n_60, n_530, n_531, n_532);
  xor g521 (n_233, A[14], A[13]);
  and g522 (n_241, A[14], A[13]);
  nand g527 (n_536, A[9], A[10]);
  xor g529 (n_537, n_233, n_210);
  xor g530 (n_237, n_537, n_235);
  nand g531 (n_538, n_233, n_210);
  nand g532 (n_539, n_235, n_210);
  nand g533 (n_540, n_233, n_235);
  nand g534 (n_245, n_538, n_539, n_540);
  xor g535 (n_541, n_236, n_237);
  xor g536 (n_26, n_541, n_238);
  nand g537 (n_542, n_236, n_237);
  nand g538 (n_543, n_238, n_237);
  nand g539 (n_544, n_236, n_238);
  nand g540 (n_59, n_542, n_543, n_544);
  xor g541 (n_240, A[15], A[14]);
  and g542 (n_246, A[15], A[14]);
  nand g547 (n_548, A[10], A[11]);
  xor g549 (n_549, n_240, n_241);
  xor g550 (n_244, n_549, n_242);
  nand g551 (n_550, n_240, n_241);
  nand g552 (n_551, n_242, n_241);
  nand g553 (n_552, n_240, n_242);
  nand g554 (n_250, n_550, n_551, n_552);
  xor g555 (n_553, n_243, n_244);
  xor g556 (n_25, n_553, n_245);
  nand g557 (n_554, n_243, n_244);
  nand g558 (n_555, n_245, n_244);
  nand g559 (n_556, n_243, n_245);
  nand g560 (n_24, n_554, n_555, n_556);
  xor g562 (n_248, n_557, A[11]);
  nand g564 (n_559, A[11], A[15]);
  nand g566 (n_251, n_558, n_559, n_560);
  xor g567 (n_561, A[12], n_246);
  xor g568 (n_249, n_561, n_247);
  nand g569 (n_562, A[12], n_246);
  nand g570 (n_563, n_247, n_246);
  nand g571 (n_564, A[12], n_247);
  nand g572 (n_253, n_562, n_563, n_564);
  xor g573 (n_565, n_248, n_249);
  xor g574 (n_58, n_565, n_250);
  nand g575 (n_566, n_248, n_249);
  nand g576 (n_567, n_250, n_249);
  nand g577 (n_568, n_248, n_250);
  nand g578 (n_23, n_566, n_567, n_568);
  xor g580 (n_252, n_169, A[12]);
  nand g582 (n_571, A[12], A[13]);
  xor g585 (n_573, n_251, n_252);
  xor g586 (n_57, n_573, n_253);
  nand g587 (n_574, n_251, n_252);
  nand g588 (n_575, n_253, n_252);
  nand g589 (n_576, n_251, n_253);
  nand g590 (n_56, n_574, n_575, n_576);
  nand g596 (n_579, n_256, n_233);
  xor g608 (n_54, n_557, n_246);
  nand g610 (n_587, n_246, A[15]);
  nand g612 (n_53, n_558, n_587, n_588);
  nand g16 (n_601, A[2], A[0]);
  xor g20 (Z[2], A[2], A[0]);
  nand g22 (n_606, A[3], A[1]);
  nand g25 (n_610, n_606, n_607, n_608);
  xor g26 (n_609, A[3], A[1]);
  nand g28 (n_611, A[4], A[2]);
  nand g29 (n_612, A[4], n_610);
  nand g30 (n_613, A[2], n_610);
  nand g31 (n_615, n_611, n_612, n_613);
  xor g32 (n_614, A[4], A[2]);
  xor g33 (Z[4], n_610, n_614);
  nand g34 (n_616, A[3], n_80);
  nand g35 (n_617, A[3], n_615);
  nand g36 (n_618, n_80, n_615);
  nand g37 (n_620, n_616, n_617, n_618);
  xor g38 (n_619, A[3], n_80);
  xor g39 (Z[5], n_615, n_619);
  nand g40 (n_621, n_45, n_79);
  nand g41 (n_622, n_45, n_620);
  nand g42 (n_623, n_79, n_620);
  nand g43 (n_625, n_621, n_622, n_623);
  xor g44 (n_624, n_45, n_79);
  xor g45 (Z[6], n_620, n_624);
  nand g46 (n_626, n_44, n_78);
  nand g47 (n_627, n_44, n_625);
  nand g48 (n_628, n_78, n_625);
  nand g49 (n_630, n_626, n_627, n_628);
  xor g50 (n_629, n_44, n_78);
  xor g51 (Z[7], n_625, n_629);
  nand g52 (n_631, n_43, n_77);
  nand g53 (n_632, n_43, n_630);
  nand g54 (n_633, n_77, n_630);
  nand g55 (n_635, n_631, n_632, n_633);
  xor g56 (n_634, n_43, n_77);
  xor g57 (Z[8], n_630, n_634);
  nand g58 (n_636, n_42, n_76);
  nand g59 (n_637, n_42, n_635);
  nand g60 (n_638, n_76, n_635);
  nand g61 (n_640, n_636, n_637, n_638);
  xor g62 (n_639, n_42, n_76);
  xor g63 (Z[9], n_635, n_639);
  nand g64 (n_641, n_41, n_75);
  nand g65 (n_642, n_41, n_640);
  nand g66 (n_643, n_75, n_640);
  nand g67 (n_645, n_641, n_642, n_643);
  xor g68 (n_644, n_41, n_75);
  xor g69 (Z[10], n_640, n_644);
  nand g70 (n_646, n_40, n_74);
  nand g71 (n_647, n_40, n_645);
  nand g72 (n_648, n_74, n_645);
  nand g73 (n_650, n_646, n_647, n_648);
  xor g74 (n_649, n_40, n_74);
  xor g75 (Z[11], n_645, n_649);
  nand g76 (n_651, n_39, n_73);
  nand g77 (n_652, n_39, n_650);
  nand g78 (n_653, n_73, n_650);
  nand g79 (n_655, n_651, n_652, n_653);
  xor g80 (n_654, n_39, n_73);
  xor g81 (Z[12], n_650, n_654);
  nand g82 (n_656, n_38, n_72);
  nand g83 (n_657, n_38, n_655);
  nand g84 (n_658, n_72, n_655);
  nand g85 (n_660, n_656, n_657, n_658);
  xor g86 (n_659, n_38, n_72);
  xor g87 (Z[13], n_655, n_659);
  nand g88 (n_661, n_37, n_71);
  nand g89 (n_662, n_37, n_660);
  nand g90 (n_663, n_71, n_660);
  nand g91 (n_665, n_661, n_662, n_663);
  xor g92 (n_664, n_37, n_71);
  xor g93 (Z[14], n_660, n_664);
  nand g94 (n_666, n_36, n_70);
  nand g95 (n_667, n_36, n_665);
  nand g96 (n_668, n_70, n_665);
  nand g97 (n_670, n_666, n_667, n_668);
  xor g618 (n_669, n_36, n_70);
  xor g619 (Z[15], n_665, n_669);
  nand g620 (n_671, n_35, n_69);
  nand g621 (n_672, n_35, n_670);
  nand g622 (n_673, n_69, n_670);
  nand g623 (n_675, n_671, n_672, n_673);
  xor g624 (n_674, n_35, n_69);
  xor g625 (Z[16], n_670, n_674);
  nand g626 (n_676, n_34, n_68);
  nand g627 (n_677, n_34, n_675);
  nand g628 (n_678, n_68, n_675);
  nand g629 (n_680, n_676, n_677, n_678);
  xor g630 (n_679, n_34, n_68);
  xor g631 (Z[17], n_675, n_679);
  nand g632 (n_681, n_33, n_67);
  nand g633 (n_682, n_33, n_680);
  nand g634 (n_683, n_67, n_680);
  nand g635 (n_685, n_681, n_682, n_683);
  xor g636 (n_684, n_33, n_67);
  xor g637 (Z[18], n_680, n_684);
  nand g638 (n_686, n_32, n_66);
  nand g639 (n_687, n_32, n_685);
  nand g640 (n_688, n_66, n_685);
  nand g641 (n_690, n_686, n_687, n_688);
  xor g642 (n_689, n_32, n_66);
  xor g643 (Z[19], n_685, n_689);
  nand g644 (n_691, n_31, n_65);
  nand g645 (n_692, n_31, n_690);
  nand g646 (n_693, n_65, n_690);
  nand g647 (n_695, n_691, n_692, n_693);
  xor g648 (n_694, n_31, n_65);
  xor g649 (Z[20], n_690, n_694);
  nand g650 (n_696, n_30, n_64);
  nand g651 (n_697, n_30, n_695);
  nand g652 (n_698, n_64, n_695);
  nand g653 (n_700, n_696, n_697, n_698);
  xor g654 (n_699, n_30, n_64);
  xor g655 (Z[21], n_695, n_699);
  nand g656 (n_701, n_29, n_63);
  nand g657 (n_702, n_29, n_700);
  nand g658 (n_703, n_63, n_700);
  nand g659 (n_705, n_701, n_702, n_703);
  xor g660 (n_704, n_29, n_63);
  xor g661 (Z[22], n_700, n_704);
  nand g662 (n_706, n_28, n_62);
  nand g663 (n_707, n_28, n_705);
  nand g664 (n_708, n_62, n_705);
  nand g665 (n_710, n_706, n_707, n_708);
  xor g666 (n_709, n_28, n_62);
  xor g667 (Z[23], n_705, n_709);
  nand g668 (n_711, n_27, n_61);
  nand g669 (n_712, n_27, n_710);
  nand g670 (n_713, n_61, n_710);
  nand g671 (n_715, n_711, n_712, n_713);
  xor g672 (n_714, n_27, n_61);
  xor g673 (Z[24], n_710, n_714);
  nand g674 (n_716, n_26, n_60);
  nand g675 (n_717, n_26, n_715);
  nand g676 (n_718, n_60, n_715);
  nand g677 (n_720, n_716, n_717, n_718);
  xor g678 (n_719, n_26, n_60);
  xor g679 (Z[25], n_715, n_719);
  nand g680 (n_721, n_25, n_59);
  nand g681 (n_722, n_25, n_720);
  nand g682 (n_723, n_59, n_720);
  nand g683 (n_725, n_721, n_722, n_723);
  xor g684 (n_724, n_25, n_59);
  xor g685 (Z[26], n_720, n_724);
  nand g686 (n_726, n_24, n_58);
  nand g687 (n_727, n_24, n_725);
  nand g688 (n_728, n_58, n_725);
  nand g689 (n_730, n_726, n_727, n_728);
  xor g690 (n_729, n_24, n_58);
  xor g691 (Z[27], n_725, n_729);
  nand g692 (n_731, n_23, n_57);
  nand g693 (n_732, n_23, n_730);
  nand g694 (n_733, n_57, n_730);
  nand g695 (n_735, n_731, n_732, n_733);
  xor g696 (n_734, n_23, n_57);
  xor g697 (Z[28], n_730, n_734);
  nand g698 (n_736, n_22, n_56);
  nand g699 (n_737, n_22, n_735);
  nand g700 (n_738, n_56, n_735);
  nand g701 (n_740, n_736, n_737, n_738);
  xor g702 (n_739, n_22, n_56);
  xor g703 (Z[29], n_735, n_739);
  nand g705 (n_742, n_21, n_740);
  nand g707 (n_745, n_741, n_742, n_743);
  xor g709 (Z[30], n_740, n_744);
  nand g710 (n_746, n_20, n_54);
  nand g711 (n_747, n_20, n_745);
  nand g712 (n_748, n_54, n_745);
  nand g713 (n_750, n_746, n_747, n_748);
  xor g714 (n_749, n_20, n_54);
  xor g715 (Z[31], n_745, n_749);
  nand g718 (n_753, n_53, n_750);
  nand g719 (n_755, n_751, n_752, n_753);
  xor g721 (Z[32], n_750, n_754);
  xnor g733 (n_357, A[16], A[14]);
  or g734 (n_358, wc, A[16]);
  not gc (wc, A[14]);
  or g735 (n_360, wc0, A[16]);
  not gc0 (wc0, A[8]);
  or g737 (n_160, n_45, A[5], A[0]);
  xnor g738 (n_163, A[9], A[5]);
  or g739 (n_170, A[5], A[9], wc1);
  not gc1 (wc1, n_387);
  xnor g740 (n_169, A[16], A[13]);
  and g741 (n_178, A[13], wc2);
  not gc2 (wc2, A[16]);
  xnor g742 (n_181, n_83, A[3]);
  xnor g744 (n_192, n_188, A[4]);
  or g747 (n_468, wc3, A[16]);
  not gc3 (wc3, A[9]);
  xnor g749 (n_229, n_382, n_521);
  or g750 (n_523, wc4, n_382);
  not gc4 (wc4, A[12]);
  or g751 (n_524, wc5, n_382);
  not gc5 (wc5, A[8]);
  xnor g752 (n_235, A[10], A[9]);
  or g753 (n_242, A[9], A[10], wc6);
  not gc6 (wc6, n_536);
  xnor g754 (n_243, A[11], A[10]);
  or g755 (n_247, A[10], A[11], wc7);
  not gc7 (wc7, n_548);
  xnor g756 (n_557, A[16], A[15]);
  or g757 (n_558, wc8, A[16]);
  not gc8 (wc8, A[15]);
  or g758 (n_560, wc9, A[16]);
  not gc9 (wc9, A[11]);
  or g759 (n_572, wc10, A[16]);
  not gc10 (wc10, A[12]);
  or g763 (n_588, A[16], wc11);
  not gc11 (wc11, n_246);
  or g764 (n_371, wc12, n_80);
  not gc12 (wc12, n_150);
  or g765 (n_372, wc13, n_80);
  not gc13 (wc13, n_149);
  or g766 (n_193, A[3], wc14, n_83);
  not gc14 (wc14, n_432);
  or g767 (n_202, A[4], wc15, n_188);
  not gc15 (wc15, n_452);
  or g768 (n_210, wc16, n_178, wc17);
  not gc17 (wc17, n_467);
  not gc16 (wc16, n_468);
  xnor g769 (n_473, n_382, n_199);
  or g770 (n_474, wc18, n_382);
  not gc18 (wc18, n_199);
  or g771 (n_476, wc19, n_382);
  not gc19 (wc19, n_200);
  xnor g772 (n_212, n_83, n_209);
  xnor g774 (n_221, n_188, n_189);
  or g775 (n_228, wc20, n_189, n_188);
  not gc20 (wc20, n_507);
  or g776 (n_256, wc21, n_178, wc22);
  not gc22 (wc22, n_571);
  not gc21 (wc21, n_572);
  or g778 (n_20, wc23, n_240, n_241);
  not gc23 (wc23, n_550);
  xnor g779 (n_156, n_80, n_369);
  or g780 (n_222, wc24, n_209, n_83);
  not gc24 (wc24, n_491);
  xnor g781 (n_22, n_233, n_256);
  or g783 (n_751, A[16], wc25);
  not gc25 (wc25, n_53);
  xnor g784 (n_754, n_53, A[16]);
  or g785 (n_21, n_256, wc26, n_233);
  not gc26 (wc26, n_579);
  or g787 (n_741, wc27, n_549);
  not gc27 (wc27, n_21);
  xnor g788 (n_744, n_549, n_21);
  or g789 (n_607, wc28, n_601);
  not gc28 (wc28, A[3]);
  or g790 (n_608, wc29, n_601);
  not gc29 (wc29, A[1]);
  xnor g791 (Z[3], n_601, n_609);
  or g792 (n_743, wc30, n_549);
  not gc30 (wc30, n_740);
  or g793 (n_752, A[16], wc31);
  not gc31 (wc31, n_750);
  not g794 (Z[33], n_755);
endmodule

module mult_signed_const_403_GENERIC(A, Z);
  input [16:0] A;
  output [33:0] Z;
  wire [16:0] A;
  wire [33:0] Z;
  mult_signed_const_403_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_527_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * -418965;"
  input [16:0] A;
  output [36:0] Z;
  wire [16:0] A;
  wire [36:0] Z;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_54, n_57;
  wire n_58, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_135, n_137;
  wire n_138, n_140, n_141, n_144, n_145, n_148, n_149, n_150;
  wire n_151, n_153, n_154, n_155, n_156, n_159, n_160, n_161;
  wire n_162, n_163, n_165, n_166, n_167, n_168, n_169, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_188, n_189, n_190, n_191;
  wire n_193, n_194, n_195, n_196, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_250, n_251, n_252, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_310, n_312, n_313;
  wire n_314, n_315, n_317, n_319, n_320, n_321, n_322, n_324;
  wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_340, n_347, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_383, n_384, n_387;
  wire n_389, n_390, n_391, n_392, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_419, n_420, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_479, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_496, n_497, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_519, n_520, n_521;
  wire n_522, n_524, n_527, n_528, n_529, n_530, n_531, n_532;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_567, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_587, n_588, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_608, n_612, n_613, n_614, n_615;
  wire n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623;
  wire n_624, n_627, n_629, n_631, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_651, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_663, n_667, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_696, n_697, n_698, n_699, n_700, n_701;
  wire n_702, n_703, n_704, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_731, n_732, n_733, n_734, n_735, n_736, n_739, n_747;
  wire n_748, n_761, n_762, n_763, n_764, n_765, n_766, n_767;
  wire n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775;
  wire n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783;
  wire n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791;
  wire n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799;
  wire n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807;
  wire n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815;
  wire n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823;
  wire n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831;
  wire n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839;
  wire n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863;
  wire n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871;
  wire n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879;
  wire n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887;
  wire n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895;
  wire n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903;
  wire n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911;
  wire n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_925;
  assign Z[0] = A[0];
  assign Z[35] = Z[36];
  xor g149 (n_87, A[0], n_135);
  xor g157 (n_86, n_349, n_138);
  nand g159 (n_351, n_138, n_137);
  nand g161 (n_48, n_350, n_351, n_352);
  xor g165 (n_85, n_353, n_141);
  nand g167 (n_355, n_141, n_140);
  nand g169 (n_47, n_354, n_355, n_356);
  nand g177 (n_150, A[0], A[3], n_360);
  xor g178 (n_361, n_144, n_145);
  nand g180 (n_362, n_144, n_145);
  nand g183 (n_46, n_362, n_363, n_364);
  xor g187 (n_151, n_365, n_148);
  nand g191 (n_156, n_366, n_367, n_368);
  xor g192 (n_369, n_149, n_150);
  xor g193 (n_83, n_369, n_151);
  nand g194 (n_370, n_149, n_150);
  nand g195 (n_371, n_151, n_150);
  nand g196 (n_372, n_149, n_151);
  nand g197 (n_45, n_370, n_371, n_372);
  xor g201 (n_155, n_373, n_153);
  nand g205 (n_162, n_374, n_375, n_376);
  xor g206 (n_377, n_154, n_155);
  xor g207 (n_82, n_377, n_156);
  nand g208 (n_378, n_154, n_155);
  nand g209 (n_379, n_156, n_155);
  nand g210 (n_380, n_154, n_156);
  nand g211 (n_44, n_378, n_379, n_380);
  nand g219 (n_166, n_360, n_383, n_384);
  nand g223 (n_387, n_160, n_159);
  xor g226 (n_389, n_161, n_162);
  xor g227 (n_81, n_389, n_163);
  nand g228 (n_390, n_161, n_162);
  nand g229 (n_391, n_163, n_162);
  nand g230 (n_392, n_161, n_163);
  nand g231 (n_43, n_390, n_391, n_392);
  nand g239 (n_173, n_366, n_395, n_396);
  xor g240 (n_397, n_54, n_165);
  xor g241 (n_169, n_397, n_166);
  nand g242 (n_398, n_54, n_165);
  nand g243 (n_399, n_166, n_165);
  nand g244 (n_400, n_54, n_166);
  nand g245 (n_176, n_398, n_399, n_400);
  xor g246 (n_401, n_167, n_168);
  xor g247 (n_80, n_401, n_169);
  nand g248 (n_402, n_167, n_168);
  nand g249 (n_403, n_169, n_168);
  nand g250 (n_404, n_167, n_169);
  nand g251 (n_42, n_402, n_403, n_404);
  nand g259 (n_181, n_374, n_407, n_408);
  xor g260 (n_409, n_171, n_172);
  xor g261 (n_175, n_409, n_173);
  nand g262 (n_410, n_171, n_172);
  nand g263 (n_411, n_173, n_172);
  nand g264 (n_412, n_171, n_173);
  nand g265 (n_184, n_410, n_411, n_412);
  xor g266 (n_413, n_174, n_175);
  xor g267 (n_79, n_413, n_176);
  nand g268 (n_414, n_174, n_175);
  nand g269 (n_415, n_176, n_175);
  nand g270 (n_416, n_174, n_176);
  nand g271 (n_41, n_414, n_415, n_416);
  nand g279 (n_190, n_384, n_419, n_420);
  xor g281 (n_183, A[0], n_179);
  xor g286 (n_425, n_180, n_181);
  xor g287 (n_185, n_425, n_182);
  nand g288 (n_426, n_180, n_181);
  nand g289 (n_427, n_182, n_181);
  nand g290 (n_428, n_180, n_182);
  nand g291 (n_195, n_426, n_427, n_428);
  xor g292 (n_429, n_183, n_184);
  xor g293 (n_78, n_429, n_185);
  nand g294 (n_430, n_183, n_184);
  nand g295 (n_431, n_185, n_184);
  nand g296 (n_432, n_183, n_185);
  nand g297 (n_40, n_430, n_431, n_432);
  nand g305 (n_200, A[7], A[4], n_396);
  nand g311 (n_201, n_438, n_439, n_440);
  xor g312 (n_441, n_188, n_189);
  xor g313 (n_194, n_441, n_190);
  nand g314 (n_442, n_188, n_189);
  nand g315 (n_443, n_190, n_189);
  nand g316 (n_444, n_188, n_190);
  nand g317 (n_204, n_442, n_443, n_444);
  xor g319 (n_196, n_445, n_193);
  nand g322 (n_448, n_191, n_193);
  nand g323 (n_206, n_446, n_447, n_448);
  xor g324 (n_449, n_194, n_195);
  xor g325 (n_77, n_449, n_196);
  nand g326 (n_450, n_194, n_195);
  nand g327 (n_451, n_196, n_195);
  nand g328 (n_452, n_194, n_196);
  nand g329 (n_39, n_450, n_451, n_452);
  nand g337 (n_210, n_408, n_455, n_456);
  xor g339 (n_203, n_457, n_198);
  nand g343 (n_214, n_458, n_459, n_460);
  xor g344 (n_461, n_199, n_200);
  xor g345 (n_205, n_461, n_201);
  nand g346 (n_462, n_199, n_200);
  nand g347 (n_463, n_201, n_200);
  nand g348 (n_464, n_199, n_201);
  nand g349 (n_215, n_462, n_463, n_464);
  xor g350 (n_465, n_202, n_203);
  xor g351 (n_207, n_465, n_204);
  nand g352 (n_466, n_202, n_203);
  nand g353 (n_467, n_204, n_203);
  nand g354 (n_468, n_202, n_204);
  nand g355 (n_218, n_466, n_467, n_468);
  xor g356 (n_469, n_205, n_206);
  xor g357 (n_76, n_469, n_207);
  nand g358 (n_470, n_205, n_206);
  nand g359 (n_471, n_207, n_206);
  nand g360 (n_472, n_205, n_207);
  nand g361 (n_38, n_470, n_471, n_472);
  nand g367 (n_221, n_474, n_475, n_476);
  nand g373 (n_220, A[6], n_479, A[12]);
  xor g375 (n_213, n_481, n_209);
  nand g379 (n_224, n_482, n_483, n_484);
  xor g380 (n_485, n_210, n_211);
  xor g381 (n_216, n_485, n_212);
  nand g382 (n_486, n_210, n_211);
  nand g383 (n_487, n_212, n_211);
  nand g384 (n_488, n_210, n_212);
  nand g385 (n_225, n_486, n_487, n_488);
  xor g386 (n_489, n_213, n_214);
  xor g387 (n_217, n_489, n_215);
  nand g388 (n_490, n_213, n_214);
  nand g389 (n_491, n_215, n_214);
  nand g390 (n_492, n_213, n_215);
  nand g391 (n_227, n_490, n_491, n_492);
  xor g392 (n_493, n_216, n_217);
  xor g393 (n_75, n_493, n_218);
  nand g394 (n_494, n_216, n_217);
  nand g395 (n_495, n_218, n_217);
  nand g396 (n_496, n_216, n_218);
  nand g397 (n_37, n_494, n_495, n_496);
  nand g405 (n_230, n_396, n_499, n_500);
  xor g407 (n_223, n_381, n_198);
  nand g411 (n_234, n_360, n_503, n_504);
  xor g412 (n_505, n_220, n_221);
  xor g413 (n_226, n_505, n_222);
  nand g414 (n_506, n_220, n_221);
  nand g415 (n_507, n_222, n_221);
  nand g416 (n_508, n_220, n_222);
  nand g417 (n_235, n_506, n_507, n_508);
  xor g418 (n_509, n_223, n_224);
  xor g419 (n_228, n_509, n_225);
  nand g420 (n_510, n_223, n_224);
  nand g421 (n_511, n_225, n_224);
  nand g422 (n_512, n_223, n_225);
  nand g423 (n_238, n_510, n_511, n_512);
  xor g424 (n_513, n_226, n_227);
  xor g425 (n_74, n_513, n_228);
  nand g426 (n_514, n_226, n_227);
  nand g427 (n_515, n_228, n_227);
  nand g428 (n_516, n_226, n_228);
  nand g429 (n_36, n_514, n_515, n_516);
  nand g435 (n_241, n_474, n_519, n_520);
  nand g441 (n_240, n_522, n_455, n_524);
  xor g443 (n_233, n_365, n_209);
  nand g447 (n_244, n_366, n_527, n_528);
  xor g448 (n_529, n_230, n_231);
  xor g449 (n_236, n_529, n_232);
  nand g450 (n_530, n_230, n_231);
  nand g451 (n_531, n_232, n_231);
  nand g452 (n_532, n_230, n_232);
  nand g453 (n_245, n_530, n_531, n_532);
  xor g454 (n_533, n_233, n_234);
  xor g455 (n_237, n_533, n_235);
  nand g456 (n_534, n_233, n_234);
  nand g457 (n_535, n_235, n_234);
  nand g458 (n_536, n_233, n_235);
  nand g459 (n_248, n_534, n_535, n_536);
  xor g460 (n_537, n_236, n_237);
  xor g461 (n_73, n_537, n_238);
  nand g462 (n_538, n_236, n_237);
  nand g463 (n_539, n_238, n_237);
  nand g464 (n_540, n_236, n_238);
  nand g465 (n_35, n_538, n_539, n_540);
  nand g473 (n_251, n_542, n_543, n_420);
  xor g475 (n_243, n_457, n_239);
  nand g479 (n_255, n_458, n_547, n_548);
  xor g480 (n_549, n_240, n_241);
  xor g481 (n_246, n_549, n_242);
  nand g482 (n_550, n_240, n_241);
  nand g483 (n_551, n_242, n_241);
  nand g484 (n_552, n_240, n_242);
  nand g485 (n_256, n_550, n_551, n_552);
  xor g486 (n_553, n_243, n_244);
  xor g487 (n_247, n_553, n_245);
  nand g488 (n_554, n_243, n_244);
  nand g489 (n_555, n_245, n_244);
  nand g490 (n_556, n_243, n_245);
  nand g491 (n_259, n_554, n_555, n_556);
  xor g492 (n_557, n_246, n_247);
  xor g493 (n_72, n_557, n_248);
  nand g494 (n_558, n_246, n_247);
  nand g495 (n_559, n_248, n_247);
  nand g496 (n_560, n_246, n_248);
  nand g497 (n_34, n_558, n_559, n_560);
  nand g503 (n_263, n_562, n_563, n_564);
  nand g509 (n_262, A[6], n_567, A[10]);
  xor g511 (n_254, n_481, n_250);
  nand g515 (n_266, n_482, n_571, n_572);
  xor g516 (n_573, n_251, n_252);
  nand g518 (n_574, n_251, n_252);
  nand g521 (n_267, n_574, n_575, n_576);
  xor g522 (n_577, n_254, n_255);
  xor g523 (n_258, n_577, n_256);
  nand g524 (n_578, n_254, n_255);
  nand g525 (n_579, n_256, n_255);
  nand g526 (n_580, n_254, n_256);
  nand g527 (n_270, n_578, n_579, n_580);
  xor g528 (n_581, n_257, n_258);
  xor g529 (n_71, n_581, n_259);
  nand g530 (n_582, n_257, n_258);
  nand g531 (n_583, n_259, n_258);
  nand g532 (n_584, n_257, n_259);
  nand g533 (n_33, n_582, n_583, n_584);
  nand g541 (n_274, n_396, n_587, n_588);
  xor g543 (n_265, A[3], n_261);
  xor g548 (n_593, n_262, n_263);
  xor g549 (n_268, n_593, n_264);
  nand g550 (n_594, n_262, n_263);
  nand g551 (n_595, n_264, n_263);
  nand g552 (n_596, n_262, n_264);
  nand g553 (n_278, n_594, n_595, n_596);
  xor g554 (n_597, n_265, n_266);
  xor g555 (n_269, n_597, n_267);
  nand g556 (n_598, n_265, n_266);
  nand g557 (n_599, n_267, n_266);
  nand g558 (n_600, n_265, n_267);
  nand g559 (n_281, n_598, n_599, n_600);
  xor g560 (n_601, n_268, n_269);
  xor g561 (n_70, n_601, n_270);
  nand g562 (n_602, n_268, n_269);
  nand g563 (n_603, n_270, n_269);
  nand g564 (n_604, n_268, n_270);
  nand g565 (n_32, n_602, n_603, n_604);
  nand g573 (n_283, n_408, n_543, n_608);
  xor g575 (n_276, A[4], n_239);
  xor g580 (n_613, n_273, n_274);
  xor g581 (n_279, n_613, n_275);
  nand g582 (n_614, n_273, n_274);
  nand g583 (n_615, n_275, n_274);
  nand g584 (n_616, n_273, n_275);
  nand g585 (n_288, n_614, n_615, n_616);
  xor g586 (n_617, n_276, n_277);
  xor g587 (n_280, n_617, n_278);
  nand g588 (n_618, n_276, n_277);
  nand g589 (n_619, n_278, n_277);
  nand g590 (n_620, n_276, n_278);
  nand g591 (n_290, n_618, n_619, n_620);
  xor g592 (n_621, n_279, n_280);
  xor g593 (n_69, n_621, n_281);
  nand g594 (n_622, n_279, n_280);
  nand g595 (n_623, n_281, n_280);
  nand g596 (n_624, n_279, n_281);
  nand g597 (n_31, n_622, n_623, n_624);
  nand g603 (n_294, n_562, n_627, n_476);
  nand g609 (n_293, n_567, n_631, n_542);
  xor g610 (n_633, n_250, n_283);
  xor g611 (n_287, n_633, n_284);
  nand g612 (n_634, n_250, n_283);
  nand g613 (n_635, n_284, n_283);
  nand g614 (n_636, n_250, n_284);
  nand g615 (n_297, n_634, n_635, n_636);
  xor g616 (n_637, n_285, n_286);
  xor g617 (n_289, n_637, n_287);
  nand g618 (n_638, n_285, n_286);
  nand g619 (n_639, n_287, n_286);
  nand g620 (n_640, n_285, n_287);
  nand g621 (n_299, n_638, n_639, n_640);
  xor g622 (n_641, n_288, n_289);
  xor g623 (n_68, n_641, n_290);
  nand g624 (n_642, n_288, n_289);
  nand g625 (n_643, n_290, n_289);
  nand g626 (n_644, n_288, n_290);
  nand g627 (n_30, n_642, n_643, n_644);
  nand g635 (n_303, n_646, n_567, n_500);
  nand g639 (n_651, n_293, n_261);
  xor g642 (n_653, n_294, n_295);
  xor g643 (n_298, n_653, n_296);
  nand g644 (n_654, n_294, n_295);
  nand g645 (n_655, n_296, n_295);
  nand g646 (n_656, n_294, n_296);
  nand g647 (n_308, n_654, n_655, n_656);
  xor g648 (n_657, n_297, n_298);
  xor g649 (n_67, n_657, n_299);
  nand g650 (n_658, n_297, n_298);
  nand g651 (n_659, n_299, n_298);
  nand g652 (n_660, n_297, n_299);
  nand g653 (n_29, n_658, n_659, n_660);
  nand g661 (n_310, n_588, n_663, n_456);
  nand g665 (n_667, n_273, n_239);
  xor g668 (n_669, n_303, n_304);
  xor g669 (n_307, n_669, n_305);
  nand g670 (n_670, n_303, n_304);
  nand g671 (n_671, n_305, n_304);
  nand g672 (n_672, n_303, n_305);
  nand g673 (n_315, n_670, n_671, n_672);
  xor g674 (n_673, n_306, n_307);
  xor g675 (n_66, n_673, n_308);
  nand g676 (n_674, n_306, n_307);
  nand g677 (n_675, n_308, n_307);
  nand g678 (n_676, n_306, n_308);
  nand g679 (n_28, n_674, n_675, n_676);
  xor g687 (n_313, n_681, n_250);
  nand g691 (n_320, n_682, n_683, n_684);
  xor g692 (n_685, n_310, n_285);
  xor g693 (n_314, n_685, n_312);
  nand g694 (n_686, n_310, n_285);
  nand g695 (n_687, n_312, n_285);
  nand g696 (n_688, n_310, n_312);
  nand g697 (n_322, n_686, n_687, n_688);
  xor g698 (n_689, n_313, n_314);
  xor g699 (n_65, n_689, n_315);
  nand g700 (n_690, n_313, n_314);
  nand g701 (n_691, n_315, n_314);
  nand g702 (n_692, n_313, n_315);
  nand g703 (n_64, n_690, n_691, n_692);
  nand g711 (n_326, A[9], A[10], n_696);
  xor g712 (n_697, n_317, n_294);
  xor g713 (n_321, n_697, n_319);
  nand g714 (n_698, n_317, n_294);
  nand g715 (n_699, n_319, n_294);
  nand g716 (n_700, n_317, n_319);
  nand g717 (n_329, n_698, n_699, n_700);
  xor g718 (n_701, n_320, n_321);
  xor g719 (n_27, n_701, n_322);
  nand g720 (n_702, n_320, n_321);
  nand g721 (n_703, n_322, n_321);
  nand g722 (n_704, n_320, n_322);
  nand g723 (n_63, n_702, n_703, n_704);
  nand g731 (n_331, A[10], A[11], n_708);
  xor g732 (n_709, n_324, n_325);
  xor g733 (n_328, n_709, n_326);
  nand g734 (n_710, n_324, n_325);
  nand g735 (n_711, n_326, n_325);
  nand g736 (n_712, n_324, n_326);
  nand g737 (n_334, n_710, n_711, n_712);
  xor g738 (n_713, n_327, n_328);
  xor g739 (n_26, n_713, n_329);
  nand g740 (n_714, n_327, n_328);
  nand g741 (n_715, n_329, n_328);
  nand g742 (n_716, n_327, n_329);
  nand g743 (n_25, n_714, n_715, n_716);
  nand g749 (n_335, n_718, n_719, n_720);
  xor g751 (n_333, n_721, n_331);
  nand g753 (n_723, n_331, n_330);
  nand g755 (n_337, n_722, n_723, n_724);
  xor g756 (n_725, n_332, n_333);
  xor g757 (n_62, n_725, n_334);
  nand g758 (n_726, n_332, n_333);
  nand g759 (n_727, n_334, n_333);
  nand g760 (n_728, n_332, n_334);
  nand g761 (n_24, n_726, n_727, n_728);
  nand g767 (n_340, n_562, n_731, n_732);
  xor g768 (n_733, n_335, n_336);
  xor g769 (n_61, n_733, n_337);
  nand g770 (n_734, n_335, n_336);
  nand g771 (n_735, n_337, n_336);
  nand g772 (n_736, n_335, n_337);
  nand g773 (n_60, n_734, n_735, n_736);
  nand g779 (n_739, n_340, n_317);
  xor g791 (n_58, n_717, n_330);
  nand g794 (n_748, A[16], n_330);
  nand g795 (n_57, n_718, n_747, n_748);
  nand g19 (n_765, n_761, n_762, n_763);
  nand g24 (n_768, n_88, n_765);
  nand g25 (n_770, n_766, n_767, n_768);
  xor g27 (Z[3], n_765, n_769);
  nand g28 (n_771, n_50, n_87);
  nand g29 (n_772, n_50, n_770);
  nand g30 (n_773, n_87, n_770);
  nand g31 (n_775, n_771, n_772, n_773);
  xor g32 (n_774, n_50, n_87);
  xor g33 (Z[4], n_770, n_774);
  nand g34 (n_776, n_49, n_86);
  nand g35 (n_777, n_49, n_775);
  nand g36 (n_778, n_86, n_775);
  nand g37 (n_780, n_776, n_777, n_778);
  xor g38 (n_779, n_49, n_86);
  xor g39 (Z[5], n_775, n_779);
  nand g40 (n_781, n_48, n_85);
  nand g41 (n_782, n_48, n_780);
  nand g42 (n_783, n_85, n_780);
  nand g43 (n_785, n_781, n_782, n_783);
  xor g44 (n_784, n_48, n_85);
  xor g45 (Z[6], n_780, n_784);
  nand g46 (n_786, n_47, n_84);
  nand g47 (n_787, n_47, n_785);
  nand g48 (n_788, n_84, n_785);
  nand g49 (n_790, n_786, n_787, n_788);
  xor g50 (n_789, n_47, n_84);
  xor g51 (Z[7], n_785, n_789);
  nand g52 (n_791, n_46, n_83);
  nand g53 (n_792, n_46, n_790);
  nand g54 (n_793, n_83, n_790);
  nand g55 (n_795, n_791, n_792, n_793);
  xor g56 (n_794, n_46, n_83);
  xor g57 (Z[8], n_790, n_794);
  nand g58 (n_796, n_45, n_82);
  nand g59 (n_797, n_45, n_795);
  nand g60 (n_798, n_82, n_795);
  nand g61 (n_800, n_796, n_797, n_798);
  xor g62 (n_799, n_45, n_82);
  xor g63 (Z[9], n_795, n_799);
  nand g64 (n_801, n_44, n_81);
  nand g65 (n_802, n_44, n_800);
  nand g66 (n_803, n_81, n_800);
  nand g67 (n_805, n_801, n_802, n_803);
  xor g68 (n_804, n_44, n_81);
  xor g69 (Z[10], n_800, n_804);
  nand g70 (n_806, n_43, n_80);
  nand g71 (n_807, n_43, n_805);
  nand g72 (n_808, n_80, n_805);
  nand g73 (n_810, n_806, n_807, n_808);
  xor g74 (n_809, n_43, n_80);
  xor g75 (Z[11], n_805, n_809);
  nand g76 (n_811, n_42, n_79);
  nand g77 (n_812, n_42, n_810);
  nand g78 (n_813, n_79, n_810);
  nand g79 (n_815, n_811, n_812, n_813);
  xor g80 (n_814, n_42, n_79);
  xor g81 (Z[12], n_810, n_814);
  nand g82 (n_816, n_41, n_78);
  nand g83 (n_817, n_41, n_815);
  nand g84 (n_818, n_78, n_815);
  nand g85 (n_820, n_816, n_817, n_818);
  xor g86 (n_819, n_41, n_78);
  xor g87 (Z[13], n_815, n_819);
  nand g88 (n_821, n_40, n_77);
  nand g89 (n_822, n_40, n_820);
  nand g90 (n_823, n_77, n_820);
  nand g91 (n_825, n_821, n_822, n_823);
  xor g92 (n_824, n_40, n_77);
  xor g93 (Z[14], n_820, n_824);
  nand g94 (n_826, n_39, n_76);
  nand g95 (n_827, n_39, n_825);
  nand g96 (n_828, n_76, n_825);
  nand g97 (n_830, n_826, n_827, n_828);
  xor g98 (n_829, n_39, n_76);
  xor g99 (Z[15], n_825, n_829);
  nand g100 (n_831, n_38, n_75);
  nand g101 (n_832, n_38, n_830);
  nand g102 (n_833, n_75, n_830);
  nand g103 (n_835, n_831, n_832, n_833);
  xor g104 (n_834, n_38, n_75);
  xor g105 (Z[16], n_830, n_834);
  nand g106 (n_836, n_37, n_74);
  nand g107 (n_837, n_37, n_835);
  nand g108 (n_838, n_74, n_835);
  nand g109 (n_840, n_836, n_837, n_838);
  xor g110 (n_839, n_37, n_74);
  xor g111 (Z[17], n_835, n_839);
  nand g112 (n_841, n_36, n_73);
  nand g113 (n_842, n_36, n_840);
  nand g114 (n_843, n_73, n_840);
  nand g115 (n_845, n_841, n_842, n_843);
  xor g116 (n_844, n_36, n_73);
  xor g117 (Z[18], n_840, n_844);
  nand g118 (n_846, n_35, n_72);
  nand g119 (n_847, n_35, n_845);
  nand g120 (n_848, n_72, n_845);
  nand g121 (n_850, n_846, n_847, n_848);
  xor g122 (n_849, n_35, n_72);
  xor g123 (Z[19], n_845, n_849);
  nand g124 (n_851, n_34, n_71);
  nand g125 (n_852, n_34, n_850);
  nand g126 (n_853, n_71, n_850);
  nand g127 (n_855, n_851, n_852, n_853);
  xor g128 (n_854, n_34, n_71);
  xor g129 (Z[20], n_850, n_854);
  nand g130 (n_856, n_33, n_70);
  nand g131 (n_857, n_33, n_855);
  nand g132 (n_858, n_70, n_855);
  nand g133 (n_860, n_856, n_857, n_858);
  xor g134 (n_859, n_33, n_70);
  xor g135 (Z[21], n_855, n_859);
  nand g136 (n_861, n_32, n_69);
  nand g137 (n_862, n_32, n_860);
  nand g138 (n_863, n_69, n_860);
  nand g139 (n_865, n_861, n_862, n_863);
  xor g140 (n_864, n_32, n_69);
  xor g141 (Z[22], n_860, n_864);
  nand g811 (n_866, n_31, n_68);
  nand g812 (n_867, n_31, n_865);
  nand g813 (n_868, n_68, n_865);
  nand g814 (n_870, n_866, n_867, n_868);
  xor g815 (n_869, n_31, n_68);
  xor g816 (Z[23], n_865, n_869);
  nand g817 (n_871, n_30, n_67);
  nand g818 (n_872, n_30, n_870);
  nand g819 (n_873, n_67, n_870);
  nand g820 (n_875, n_871, n_872, n_873);
  xor g821 (n_874, n_30, n_67);
  xor g822 (Z[24], n_870, n_874);
  nand g823 (n_876, n_29, n_66);
  nand g824 (n_877, n_29, n_875);
  nand g825 (n_878, n_66, n_875);
  nand g826 (n_880, n_876, n_877, n_878);
  xor g827 (n_879, n_29, n_66);
  xor g828 (Z[25], n_875, n_879);
  nand g829 (n_881, n_28, n_65);
  nand g830 (n_882, n_28, n_880);
  nand g831 (n_883, n_65, n_880);
  nand g832 (n_885, n_881, n_882, n_883);
  xor g833 (n_884, n_28, n_65);
  xor g834 (Z[26], n_880, n_884);
  nand g835 (n_886, n_27, n_64);
  nand g836 (n_887, n_27, n_885);
  nand g837 (n_888, n_64, n_885);
  nand g838 (n_890, n_886, n_887, n_888);
  xor g839 (n_889, n_27, n_64);
  xor g840 (Z[27], n_885, n_889);
  nand g841 (n_891, n_26, n_63);
  nand g842 (n_892, n_26, n_890);
  nand g843 (n_893, n_63, n_890);
  nand g844 (n_895, n_891, n_892, n_893);
  xor g845 (n_894, n_26, n_63);
  xor g846 (Z[28], n_890, n_894);
  nand g847 (n_896, n_25, n_62);
  nand g848 (n_897, n_25, n_895);
  nand g849 (n_898, n_62, n_895);
  nand g850 (n_900, n_896, n_897, n_898);
  xor g851 (n_899, n_25, n_62);
  xor g852 (Z[29], n_895, n_899);
  nand g853 (n_901, n_24, n_61);
  nand g854 (n_902, n_24, n_900);
  nand g855 (n_903, n_61, n_900);
  nand g856 (n_905, n_901, n_902, n_903);
  xor g857 (n_904, n_24, n_61);
  xor g858 (Z[30], n_900, n_904);
  nand g859 (n_906, n_23, n_60);
  nand g860 (n_907, n_23, n_905);
  nand g861 (n_908, n_60, n_905);
  nand g862 (n_910, n_906, n_907, n_908);
  xor g863 (n_909, n_23, n_60);
  xor g864 (Z[31], n_905, n_909);
  nand g866 (n_912, n_22, n_910);
  nand g868 (n_915, n_911, n_912, n_913);
  xor g870 (Z[32], n_910, n_914);
  nand g871 (n_916, n_21, n_58);
  nand g872 (n_917, n_21, n_915);
  nand g873 (n_918, n_58, n_915);
  nand g874 (n_920, n_916, n_917, n_918);
  xor g875 (n_919, n_21, n_58);
  xor g876 (Z[33], n_915, n_919);
  nand g877 (n_921, A[16], n_57);
  nand g878 (n_922, A[16], n_920);
  nand g879 (n_923, n_57, n_920);
  nand g880 (n_925, n_921, n_922, n_923);
  xor g881 (n_924, A[16], n_57);
  xor g882 (Z[34], n_920, n_924);
  xor g891 (n_88, A[3], A[1]);
  nor g892 (n_50, A[3], A[1]);
  xor g893 (n_135, A[4], A[2]);
  nor g894 (n_138, A[4], A[2]);
  xor g895 (n_137, A[5], A[3]);
  nor g896 (n_141, A[5], A[3]);
  xor g897 (n_140, A[6], A[4]);
  nor g898 (n_145, A[6], A[4]);
  xor g899 (n_144, A[7], A[5]);
  nor g900 (n_148, A[7], A[5]);
  or g901 (n_360, A[3], A[0]);
  xor g902 (n_149, A[8], A[6]);
  nor g903 (n_153, A[8], A[6]);
  xor g904 (n_365, A[4], A[1]);
  or g905 (n_366, A[4], A[1]);
  xor g906 (n_154, A[9], A[7]);
  nor g907 (n_160, A[9], A[7]);
  xor g908 (n_373, A[5], A[2]);
  or g909 (n_374, A[5], A[2]);
  xor g910 (n_159, A[10], A[8]);
  nor g911 (n_165, A[10], A[8]);
  xor g912 (n_381, A[3], A[0]);
  or g913 (n_383, A[6], A[0]);
  or g914 (n_384, A[6], A[3]);
  xor g915 (n_54, A[11], A[9]);
  nor g916 (n_172, A[11], A[9]);
  or g917 (n_395, A[7], A[1]);
  or g918 (n_396, A[7], A[4]);
  xor g919 (n_171, A[12], A[10]);
  nor g920 (n_179, A[12], A[10]);
  or g921 (n_407, A[8], A[2]);
  or g922 (n_408, A[8], A[5]);
  xor g923 (n_180, A[13], A[11]);
  nor g924 (n_188, A[13], A[11]);
  xor g925 (n_417, A[6], A[3]);
  or g926 (n_419, A[9], A[3]);
  or g927 (n_420, A[9], A[6]);
  xor g928 (n_189, A[14], A[12]);
  nor g929 (n_199, A[14], A[12]);
  xor g930 (n_437, A[10], A[1]);
  or g931 (n_438, A[10], A[1]);
  or g932 (n_439, A[1], A[0]);
  or g933 (n_440, A[10], A[0]);
  xor g934 (n_198, A[15], A[13]);
  nor g935 (n_209, A[15], A[13]);
  xor g936 (n_453, A[8], A[5]);
  or g937 (n_455, A[11], A[5]);
  or g938 (n_456, A[11], A[8]);
  xor g939 (n_457, A[2], A[1]);
  or g940 (n_458, A[2], A[1]);
  xnor g941 (n_473, A[16], A[14]);
  or g942 (n_474, A[14], wc);
  not gc (wc, A[16]);
  or g943 (n_475, A[14], A[9]);
  or g944 (n_476, A[9], wc0);
  not gc0 (wc0, A[16]);
  or g945 (n_479, A[12], A[6]);
  xor g946 (n_481, A[3], A[2]);
  or g947 (n_482, A[3], A[2]);
  xor g948 (n_497, A[7], A[4]);
  or g949 (n_499, A[10], A[4]);
  or g950 (n_500, A[10], A[7]);
  or g951 (n_519, A[14], A[8]);
  or g952 (n_520, A[8], wc1);
  not gc1 (wc1, A[16]);
  xor g953 (n_521, A[5], A[0]);
  or g954 (n_522, A[5], A[0]);
  or g955 (n_524, A[11], A[0]);
  xor g956 (n_239, A[15], A[12]);
  nor g957 (n_250, A[15], A[12]);
  xor g958 (n_541, A[6], A[5]);
  or g959 (n_542, A[6], A[5]);
  or g960 (n_543, A[9], A[5]);
  xnor g961 (n_561, A[16], A[13]);
  or g962 (n_562, A[13], wc2);
  not gc2 (wc2, A[16]);
  or g963 (n_563, A[13], A[7]);
  or g964 (n_564, A[7], wc3);
  not gc3 (wc3, A[16]);
  or g965 (n_567, A[10], A[6]);
  xor g966 (n_261, A[14], A[11]);
  nor g967 (n_273, A[14], A[11]);
  or g968 (n_587, A[8], A[4]);
  or g969 (n_588, A[8], A[7]);
  or g970 (n_608, A[9], A[8]);
  or g971 (n_627, A[13], A[9]);
  xor g972 (n_629, A[10], A[6]);
  or g973 (n_631, A[10], A[5]);
  xor g974 (n_645, A[7], A[6]);
  or g975 (n_646, A[7], A[6]);
  xor g976 (n_661, A[8], A[7]);
  or g977 (n_663, A[11], A[7]);
  xor g978 (n_681, A[12], A[8]);
  or g979 (n_682, A[12], A[8]);
  xor g980 (n_317, A[14], A[13]);
  nor g981 (n_325, A[14], A[13]);
  or g982 (n_696, A[10], A[9]);
  xor g983 (n_324, A[15], A[14]);
  nor g984 (n_330, A[15], A[14]);
  or g985 (n_708, A[11], A[10]);
  xnor g986 (n_717, A[16], A[15]);
  or g987 (n_718, A[15], wc4);
  not gc4 (wc4, A[16]);
  or g988 (n_719, A[15], A[11]);
  or g989 (n_720, A[11], wc5);
  not gc5 (wc5, A[16]);
  or g990 (n_731, A[13], A[12]);
  or g991 (n_732, A[12], wc6);
  not gc6 (wc6, A[16]);
  or g992 (n_347, A[0], wc7);
  not gc7 (wc7, n_135);
  xnor g994 (n_349, n_137, A[1]);
  or g995 (n_350, A[1], wc8);
  not gc8 (wc8, n_137);
  or g996 (n_352, A[1], wc9);
  not gc9 (wc9, n_138);
  xnor g997 (n_353, n_140, A[2]);
  or g998 (n_354, A[2], wc10);
  not gc10 (wc10, n_140);
  or g999 (n_356, A[2], wc11);
  not gc11 (wc11, n_141);
  or g1001 (n_367, A[4], wc12);
  not gc12 (wc12, n_148);
  or g1002 (n_368, A[1], wc13);
  not gc13 (wc13, n_148);
  or g1003 (n_375, A[5], wc14);
  not gc14 (wc14, n_153);
  or g1004 (n_376, A[2], wc15);
  not gc15 (wc15, n_153);
  xnor g1005 (n_161, n_381, A[6]);
  xnor g1008 (n_167, n_365, A[7]);
  xnor g1009 (n_174, n_373, A[8]);
  xnor g1010 (n_182, n_417, A[9]);
  or g1012 (n_424, A[0], wc16);
  not gc16 (wc16, n_179);
  xnor g1014 (n_191, n_437, A[0]);
  xnor g1015 (n_202, n_453, A[11]);
  or g1016 (n_459, A[1], wc17);
  not gc17 (wc17, n_198);
  or g1017 (n_460, A[2], wc18);
  not gc18 (wc18, n_198);
  xnor g1018 (n_211, n_473, A[9]);
  xnor g1019 (n_212, A[12], A[6]);
  or g1020 (n_483, A[2], wc19);
  not gc19 (wc19, n_209);
  or g1021 (n_484, A[3], wc20);
  not gc20 (wc20, n_209);
  xnor g1022 (n_222, n_497, A[10]);
  or g1023 (n_503, A[0], wc21);
  not gc21 (wc21, n_198);
  or g1024 (n_504, A[3], wc22);
  not gc22 (wc22, n_198);
  xnor g1025 (n_231, n_473, A[8]);
  xnor g1026 (n_232, n_521, A[11]);
  or g1027 (n_527, A[1], wc23);
  not gc23 (wc23, n_209);
  or g1028 (n_528, A[4], wc24);
  not gc24 (wc24, n_209);
  xnor g1029 (n_242, n_541, A[9]);
  or g1030 (n_547, A[1], wc25);
  not gc25 (wc25, n_239);
  or g1031 (n_548, A[2], wc26);
  not gc26 (wc26, n_239);
  xnor g1032 (n_252, n_561, A[7]);
  or g1034 (n_571, A[2], wc27);
  not gc27 (wc27, n_250);
  or g1035 (n_572, A[3], wc28);
  not gc28 (wc28, n_250);
  xnor g1036 (n_264, n_497, A[8]);
  or g1038 (n_592, A[3], wc29);
  not gc29 (wc29, n_261);
  xnor g1039 (n_275, n_453, A[9]);
  or g1041 (n_612, A[4], wc30);
  not gc30 (wc30, n_239);
  xnor g1042 (n_285, n_561, A[9]);
  xnor g1043 (n_284, n_629, A[5]);
  xnor g1044 (n_295, n_645, A[10]);
  xnor g1045 (n_304, n_661, A[11]);
  or g1047 (n_683, A[12], wc31);
  not gc31 (wc31, n_250);
  or g1048 (n_684, A[8], wc32);
  not gc32 (wc32, n_250);
  xnor g1049 (n_319, A[10], A[9]);
  xnor g1050 (n_327, A[11], A[10]);
  xnor g1051 (n_332, n_717, A[11]);
  xnor g1052 (n_721, n_330, A[12]);
  or g1053 (n_722, A[12], wc33);
  not gc33 (wc33, n_330);
  xnor g1054 (n_336, n_561, A[12]);
  or g1058 (n_747, A[15], wc34);
  not gc34 (wc34, n_330);
  or g1059 (n_761, A[0], wc35);
  not gc35 (wc35, A[2]);
  xnor g1060 (n_764, A[2], A[0]);
  or g1061 (n_766, A[2], wc36);
  not gc36 (wc36, n_88);
  xnor g1062 (n_769, n_88, A[2]);
  or g1063 (n_49, wc37, wc38, n_135);
  not gc38 (wc38, n_347);
  not gc37 (wc37, A[0]);
  xnor g1064 (n_84, n_361, n_381);
  or g1065 (n_363, n_381, wc39);
  not gc39 (wc39, n_145);
  or g1066 (n_364, n_381, wc40);
  not gc40 (wc40, n_144);
  xnor g1067 (n_163, n_160, n_159);
  or g1068 (n_168, n_159, n_160, wc41);
  not gc41 (wc41, n_387);
  or g1069 (n_193, wc42, wc43, n_179);
  not gc43 (wc43, n_424);
  not gc42 (wc42, A[0]);
  xnor g1070 (n_445, n_497, n_191);
  or g1071 (n_446, wc44, n_497);
  not gc44 (wc44, n_191);
  or g1072 (n_575, wc45, n_629);
  not gc45 (wc45, n_252);
  or g1073 (n_576, n_629, wc46);
  not gc46 (wc46, n_251);
  or g1074 (n_277, wc47, wc48, n_261);
  not gc48 (wc48, n_592);
  not gc47 (wc47, A[3]);
  or g1075 (n_286, wc49, wc50, n_239);
  not gc50 (wc50, n_612);
  not gc49 (wc49, A[4]);
  xnor g1076 (n_296, n_293, n_261);
  xnor g1078 (n_305, n_239, n_273);
  or g1079 (n_312, n_273, n_239, wc51);
  not gc51 (wc51, n_667);
  or g1080 (n_724, A[12], wc52);
  not gc52 (wc52, n_331);
  xnor g1081 (n_23, n_340, n_317);
  or g1084 (n_21, n_324, n_325, wc53);
  not gc53 (wc53, n_710);
  xor g1085 (Z[1], A[1], A[0]);
  or g1086 (n_447, wc54, n_497);
  not gc54 (wc54, n_193);
  xnor g1087 (n_257, n_573, n_629);
  or g1088 (n_306, n_261, wc55, n_293);
  not gc55 (wc55, n_651);
  or g1089 (n_22, n_317, wc56, n_340);
  not gc56 (wc56, n_739);
  or g1091 (n_762, n_439, A[0]);
  or g1092 (n_763, wc57, n_439);
  not gc57 (wc57, A[2]);
  xnor g1093 (Z[2], n_439, n_764);
  or g1094 (n_911, wc58, n_709);
  not gc58 (wc58, n_22);
  xnor g1095 (n_914, n_709, n_22);
  or g1096 (n_767, A[2], wc59);
  not gc59 (wc59, n_765);
  or g1097 (n_913, wc60, n_709);
  not gc60 (wc60, n_910);
  not g1098 (Z[36], n_925);
endmodule

module mult_signed_const_527_GENERIC(A, Z);
  input [16:0] A;
  output [36:0] Z;
  wire [16:0] A;
  wire [36:0] Z;
  mult_signed_const_527_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_608_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 41429;"
  input [16:0] A;
  output [32:0] Z;
  wire [16:0] A;
  wire [32:0] Z;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_45;
  wire n_47, n_48, n_49, n_50, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_81;
  wire n_120, n_122, n_123, n_125, n_126, n_128, n_129, n_130;
  wire n_132, n_133, n_134, n_135, n_137, n_138, n_139, n_140;
  wire n_142, n_143, n_144, n_145, n_146, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_213, n_214, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_225, n_226, n_227, n_228, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_239, n_241;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_333, n_334, n_335, n_336, n_337, n_338, n_340;
  wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_349, n_350, n_351, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_367, n_368;
  wire n_369, n_371, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_406, n_407, n_408;
  wire n_409, n_410, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_426, n_427;
  wire n_430, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_478, n_479, n_482, n_484, n_485, n_486;
  wire n_487, n_490, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_499, n_500, n_501, n_502, n_503, n_506, n_510, n_514;
  wire n_518, n_519, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567;
  wire n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575;
  wire n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591;
  wire n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599;
  wire n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615;
  wire n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623;
  wire n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631;
  wire n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639;
  wire n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647;
  wire n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655;
  wire n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663;
  wire n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679;
  wire n_680, n_681;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g100 (n_79, A[4], A[0]);
  and g101 (n_45, A[4], A[0]);
  xor g102 (n_248, A[5], A[3]);
  xor g103 (n_78, n_248, A[1]);
  nand g104 (n_249, A[5], A[3]);
  nand g105 (n_250, A[1], A[3]);
  nand g106 (n_251, A[5], A[1]);
  nand g107 (n_120, n_249, n_250, n_251);
  xor g108 (n_252, A[6], A[4]);
  nand g110 (n_253, A[6], A[4]);
  nand g117 (n_258, n_120, A[2]);
  nand g119 (n_43, n_257, n_258, n_259);
  xor g120 (n_260, A[7], A[5]);
  nand g122 (n_261, A[7], A[5]);
  nand g125 (n_125, n_261, n_262, n_263);
  xor g126 (n_264, A[3], n_122);
  xor g127 (n_76, n_264, n_123);
  nand g128 (n_265, A[3], n_122);
  nand g129 (n_266, n_123, n_122);
  nand g130 (n_267, A[3], n_123);
  nand g131 (n_42, n_265, n_266, n_267);
  xor g132 (n_268, A[8], A[6]);
  nand g134 (n_269, A[8], A[6]);
  nand g137 (n_129, n_269, n_270, n_271);
  xor g138 (n_272, A[4], n_125);
  xor g139 (n_75, n_272, n_126);
  nand g140 (n_273, A[4], n_125);
  nand g141 (n_274, n_126, n_125);
  nand g142 (n_275, A[4], n_126);
  nand g143 (n_41, n_273, n_274, n_275);
  xor g144 (n_128, A[9], A[7]);
  and g145 (n_132, A[9], A[7]);
  xor g147 (n_130, n_276, A[5]);
  nand g149 (n_278, A[5], A[0]);
  nand g151 (n_133, n_277, n_278, n_279);
  xor g152 (n_280, n_128, n_129);
  xor g153 (n_74, n_280, n_130);
  nand g154 (n_281, n_128, n_129);
  nand g155 (n_282, n_130, n_129);
  nand g156 (n_283, n_128, n_130);
  nand g157 (n_40, n_281, n_282, n_283);
  xor g158 (n_284, A[10], A[8]);
  nand g160 (n_285, A[10], A[8]);
  nand g163 (n_137, n_285, n_286, n_287);
  xor g164 (n_288, A[1], A[6]);
  xor g165 (n_135, n_288, n_132);
  nand g166 (n_289, A[1], A[6]);
  nand g167 (n_290, n_132, A[6]);
  nand g168 (n_291, A[1], n_132);
  nand g169 (n_139, n_289, n_290, n_291);
  xor g170 (n_292, n_133, n_134);
  xor g171 (n_73, n_292, n_135);
  nand g172 (n_293, n_133, n_134);
  nand g173 (n_294, n_135, n_134);
  nand g174 (n_295, n_133, n_135);
  nand g175 (n_39, n_293, n_294, n_295);
  xor g176 (n_296, A[11], A[9]);
  nand g178 (n_297, A[11], A[9]);
  nand g181 (n_142, n_297, n_298, n_299);
  xor g182 (n_300, A[2], A[7]);
  xor g183 (n_140, n_300, n_137);
  nand g184 (n_301, A[2], A[7]);
  nand g185 (n_302, n_137, A[7]);
  nand g186 (n_303, A[2], n_137);
  nand g187 (n_145, n_301, n_302, n_303);
  xor g188 (n_304, n_138, n_139);
  xor g189 (n_72, n_304, n_140);
  nand g190 (n_305, n_138, n_139);
  nand g191 (n_306, n_140, n_139);
  nand g192 (n_307, n_138, n_140);
  nand g193 (n_38, n_305, n_306, n_307);
  xor g194 (n_308, A[12], A[10]);
  nand g196 (n_309, A[12], A[10]);
  nand g199 (n_48, n_309, n_310, n_311);
  xor g200 (n_312, A[3], A[8]);
  xor g201 (n_144, n_312, n_142);
  nand g202 (n_313, A[3], A[8]);
  nand g203 (n_314, n_142, A[8]);
  nand g204 (n_315, A[3], n_142);
  nand g205 (n_146, n_313, n_314, n_315);
  xor g206 (n_316, n_143, n_144);
  xor g207 (n_71, n_316, n_145);
  nand g208 (n_317, n_143, n_144);
  nand g209 (n_318, n_145, n_144);
  nand g210 (n_319, n_143, n_145);
  nand g211 (n_37, n_317, n_318, n_319);
  xor g212 (n_47, A[13], A[11]);
  and g213 (n_148, A[13], A[11]);
  xor g215 (n_49, n_320, A[9]);
  nand g217 (n_322, A[9], A[4]);
  nand g219 (n_149, n_321, n_322, n_323);
  xor g220 (n_324, A[0], n_47);
  xor g221 (n_50, n_324, n_48);
  nand g222 (n_325, A[0], n_47);
  nand g223 (n_326, n_48, n_47);
  nand g224 (n_327, A[0], n_48);
  nand g225 (n_152, n_325, n_326, n_327);
  xor g226 (n_328, n_49, n_50);
  xor g227 (n_70, n_328, n_146);
  nand g228 (n_329, n_49, n_50);
  nand g229 (n_330, n_146, n_50);
  nand g230 (n_331, n_49, n_146);
  nand g231 (n_36, n_329, n_330, n_331);
  xor g232 (n_241, A[14], A[12]);
  nand g234 (n_333, A[14], A[12]);
  nand g237 (n_156, n_333, n_334, n_335);
  xor g238 (n_336, A[5], A[10]);
  xor g239 (n_151, n_336, A[1]);
  nand g240 (n_337, A[5], A[10]);
  nand g241 (n_338, A[1], A[10]);
  nand g243 (n_157, n_337, n_338, n_251);
  xor g244 (n_340, n_148, n_149);
  xor g245 (n_153, n_340, n_150);
  nand g246 (n_341, n_148, n_149);
  nand g247 (n_342, n_150, n_149);
  nand g248 (n_343, n_148, n_150);
  nand g249 (n_161, n_341, n_342, n_343);
  xor g250 (n_344, n_151, n_152);
  xor g251 (n_69, n_344, n_153);
  nand g252 (n_345, n_151, n_152);
  nand g253 (n_346, n_153, n_152);
  nand g254 (n_347, n_151, n_153);
  nand g255 (n_35, n_345, n_346, n_347);
  xor g256 (n_81, A[15], A[13]);
  and g257 (n_164, A[15], A[13]);
  xor g259 (n_158, n_348, A[11]);
  nand g261 (n_350, A[11], A[6]);
  nand g263 (n_166, n_349, n_350, n_351);
  xor g264 (Z[2], A[2], A[0]);
  xor g265 (n_159, Z[2], n_81);
  nand g266 (n_353, A[2], A[0]);
  nand g267 (n_354, n_81, A[0]);
  nand g268 (n_355, A[2], n_81);
  nand g269 (n_169, n_353, n_354, n_355);
  xor g270 (n_356, n_156, n_157);
  xor g271 (n_160, n_356, n_158);
  nand g272 (n_357, n_156, n_157);
  nand g273 (n_358, n_158, n_157);
  nand g274 (n_359, n_156, n_158);
  nand g275 (n_171, n_357, n_358, n_359);
  xor g276 (n_360, n_159, n_160);
  xor g277 (n_68, n_360, n_161);
  nand g278 (n_361, n_159, n_160);
  nand g279 (n_362, n_161, n_160);
  nand g280 (n_363, n_159, n_161);
  nand g281 (n_34, n_361, n_362, n_363);
  xor g285 (n_168, A[10], A[7]);
  xor g290 (n_368, A[12], A[3]);
  xor g291 (n_167, n_368, A[1]);
  nand g292 (n_369, A[12], A[3]);
  nand g294 (n_371, A[12], A[1]);
  nand g295 (n_176, n_369, n_250, n_371);
  xor g296 (n_54, n_164, n_165);
  xor g297 (n_170, n_54, n_166);
  nand g298 (n_373, n_164, n_165);
  nand g299 (n_374, n_166, n_165);
  nand g300 (n_375, n_164, n_166);
  nand g301 (n_179, n_373, n_374, n_375);
  xor g302 (n_376, n_167, n_168);
  xor g303 (n_172, n_376, n_169);
  nand g304 (n_377, n_167, n_168);
  nand g305 (n_378, n_169, n_168);
  nand g306 (n_379, n_167, n_169);
  nand g307 (n_181, n_377, n_378, n_379);
  xor g308 (n_380, n_170, n_171);
  xor g309 (n_67, n_380, n_172);
  nand g310 (n_381, n_170, n_171);
  nand g311 (n_382, n_172, n_171);
  nand g312 (n_383, n_170, n_172);
  nand g313 (n_33, n_381, n_382, n_383);
  xor g316 (n_384, A[8], A[4]);
  nand g318 (n_385, A[8], A[4]);
  nand g321 (n_185, n_385, n_386, n_387);
  xor g328 (n_392, n_174, n_175);
  xor g329 (n_180, n_392, n_176);
  nand g330 (n_393, n_174, n_175);
  nand g331 (n_394, n_176, n_175);
  nand g332 (n_395, n_174, n_176);
  nand g333 (n_189, n_393, n_394, n_395);
  xor g334 (n_396, n_177, n_178);
  xor g335 (n_182, n_396, n_179);
  nand g336 (n_397, n_177, n_178);
  nand g337 (n_398, n_179, n_178);
  nand g338 (n_399, n_177, n_179);
  nand g339 (n_192, n_397, n_398, n_399);
  xor g340 (n_400, n_180, n_181);
  xor g341 (n_66, n_400, n_182);
  nand g342 (n_401, n_180, n_181);
  nand g343 (n_402, n_182, n_181);
  nand g344 (n_403, n_180, n_182);
  nand g345 (n_32, n_401, n_402, n_403);
  xor g347 (n_187, n_165, A[9]);
  nand g349 (n_406, A[9], A[14]);
  xor g353 (n_186, n_408, A[3]);
  nand g357 (n_196, n_409, n_410, n_249);
  xor g358 (n_412, n_164, n_185);
  xor g359 (n_190, n_412, n_186);
  nand g360 (n_413, n_164, n_185);
  nand g361 (n_414, n_186, n_185);
  nand g362 (n_415, n_164, n_186);
  nand g363 (n_200, n_413, n_414, n_415);
  xor g364 (n_416, n_187, n_188);
  xor g365 (n_191, n_416, n_189);
  nand g366 (n_417, n_187, n_188);
  nand g367 (n_418, n_189, n_188);
  nand g368 (n_419, n_187, n_189);
  nand g369 (n_202, n_417, n_418, n_419);
  xor g370 (n_420, n_190, n_191);
  xor g371 (n_65, n_420, n_192);
  nand g372 (n_421, n_190, n_191);
  nand g373 (n_422, n_192, n_191);
  nand g374 (n_423, n_190, n_192);
  nand g375 (n_31, n_421, n_422, n_423);
  xor g379 (n_198, n_252, A[10]);
  nand g381 (n_426, A[10], A[4]);
  nand g382 (n_427, A[6], A[10]);
  nand g383 (n_205, n_253, n_426, n_427);
  xor g385 (n_199, n_81, n_196);
  xor g390 (n_432, n_197, n_198);
  xor g391 (n_201, n_432, n_199);
  nand g392 (n_433, n_197, n_198);
  nand g393 (n_434, n_199, n_198);
  nand g394 (n_435, n_197, n_199);
  nand g395 (n_210, n_433, n_434, n_435);
  xor g396 (n_436, n_200, n_201);
  xor g397 (n_64, n_436, n_202);
  nand g398 (n_437, n_200, n_201);
  nand g399 (n_438, n_202, n_201);
  nand g400 (n_439, n_200, n_202);
  nand g401 (n_30, n_437, n_438, n_439);
  nand g407 (n_214, n_441, n_442, n_443);
  xor g408 (n_444, A[5], A[11]);
  xor g409 (n_207, n_444, n_204);
  nand g410 (n_445, A[5], A[11]);
  nand g411 (n_446, n_204, A[11]);
  nand g412 (n_447, A[5], n_204);
  nand g413 (n_216, n_445, n_446, n_447);
  xor g414 (n_448, n_205, n_206);
  xor g415 (n_209, n_448, n_207);
  nand g416 (n_449, n_205, n_206);
  nand g417 (n_450, n_207, n_206);
  nand g418 (n_451, n_205, n_207);
  nand g419 (n_218, n_449, n_450, n_451);
  xor g420 (n_452, n_208, n_209);
  xor g421 (n_63, n_452, n_210);
  nand g422 (n_453, n_208, n_209);
  nand g423 (n_454, n_210, n_209);
  nand g424 (n_455, n_208, n_210);
  nand g425 (n_62, n_453, n_454, n_455);
  xor g434 (n_460, n_213, n_214);
  nand g436 (n_461, n_213, n_214);
  nand g439 (n_223, n_461, n_462, n_463);
  xor g440 (n_464, n_216, n_217);
  xor g441 (n_29, n_464, n_218);
  nand g442 (n_465, n_216, n_217);
  nand g443 (n_466, n_218, n_217);
  nand g444 (n_467, n_216, n_218);
  nand g445 (n_61, n_465, n_466, n_467);
  xor g446 (n_468, A[16], A[13]);
  xor g447 (n_221, n_468, A[7]);
  nand g448 (n_469, A[16], A[13]);
  nand g449 (n_470, A[7], A[13]);
  nand g450 (n_471, A[16], A[7]);
  nand g451 (n_226, n_469, n_470, n_471);
  xor g452 (n_472, A[9], n_219);
  xor g453 (n_222, n_472, n_220);
  nand g454 (n_473, A[9], n_219);
  nand g455 (n_474, n_220, n_219);
  nand g456 (n_475, A[9], n_220);
  nand g457 (n_228, n_473, n_474, n_475);
  xor g458 (n_476, n_221, n_222);
  xor g459 (n_28, n_476, n_223);
  nand g460 (n_477, n_221, n_222);
  nand g461 (n_478, n_223, n_222);
  nand g462 (n_479, n_221, n_223);
  nand g463 (n_60, n_477, n_478, n_479);
  xor g464 (n_225, A[14], A[10]);
  and g465 (n_230, A[14], A[10]);
  nand g469 (n_482, n_225, A[8]);
  xor g472 (n_484, n_226, n_227);
  xor g473 (n_27, n_484, n_228);
  nand g474 (n_485, n_226, n_227);
  nand g475 (n_486, n_228, n_227);
  nand g476 (n_487, n_226, n_228);
  nand g477 (n_26, n_485, n_486, n_487);
  xor g478 (n_231, A[15], A[11]);
  and g479 (n_234, A[15], A[11]);
  nand g483 (n_490, n_230, A[9]);
  xor g486 (n_492, n_231, n_232);
  xor g487 (n_59, n_492, n_233);
  nand g488 (n_493, n_231, n_232);
  nand g489 (n_494, n_233, n_232);
  nand g490 (n_495, n_231, n_233);
  nand g491 (n_25, n_493, n_494, n_495);
  xor g493 (n_235, n_496, A[10]);
  nand g497 (n_239, n_497, n_309, n_499);
  xor g498 (n_500, n_234, n_235);
  xor g499 (n_58, n_500, n_236);
  nand g500 (n_501, n_234, n_235);
  nand g501 (n_502, n_236, n_235);
  nand g502 (n_503, n_234, n_236);
  nand g503 (n_57, n_501, n_502, n_503);
  nand g509 (n_506, n_239, n_47);
  nand g517 (n_510, n_148, n_241);
  nand g531 (n_518, n_164, A[14]);
  nand g25 (n_541, n_250, n_538, n_539);
  xor g26 (n_540, A[3], A[1]);
  nand g28 (n_542, A[2], n_79);
  nand g29 (n_543, A[2], n_541);
  nand g30 (n_544, n_79, n_541);
  nand g31 (n_546, n_542, n_543, n_544);
  xor g32 (n_545, A[2], n_79);
  xor g33 (Z[4], n_541, n_545);
  nand g34 (n_547, n_45, n_78);
  nand g35 (n_548, n_45, n_546);
  nand g36 (n_549, n_78, n_546);
  nand g37 (n_551, n_547, n_548, n_549);
  xor g38 (n_550, n_45, n_78);
  xor g39 (Z[5], n_546, n_550);
  nand g42 (n_554, n_77, n_551);
  nand g43 (n_556, n_552, n_553, n_554);
  xor g45 (Z[6], n_551, n_555);
  nand g46 (n_557, n_43, n_76);
  nand g47 (n_558, n_43, n_556);
  nand g48 (n_559, n_76, n_556);
  nand g49 (n_561, n_557, n_558, n_559);
  xor g50 (n_560, n_43, n_76);
  xor g51 (Z[7], n_556, n_560);
  nand g52 (n_562, n_42, n_75);
  nand g53 (n_563, n_42, n_561);
  nand g54 (n_564, n_75, n_561);
  nand g55 (n_566, n_562, n_563, n_564);
  xor g56 (n_565, n_42, n_75);
  xor g57 (Z[8], n_561, n_565);
  nand g58 (n_567, n_41, n_74);
  nand g59 (n_568, n_41, n_566);
  nand g60 (n_569, n_74, n_566);
  nand g61 (n_571, n_567, n_568, n_569);
  xor g62 (n_570, n_41, n_74);
  xor g63 (Z[9], n_566, n_570);
  nand g64 (n_572, n_40, n_73);
  nand g65 (n_573, n_40, n_571);
  nand g66 (n_574, n_73, n_571);
  nand g67 (n_576, n_572, n_573, n_574);
  xor g68 (n_575, n_40, n_73);
  xor g69 (Z[10], n_571, n_575);
  nand g70 (n_577, n_39, n_72);
  nand g71 (n_578, n_39, n_576);
  nand g72 (n_579, n_72, n_576);
  nand g73 (n_581, n_577, n_578, n_579);
  xor g74 (n_580, n_39, n_72);
  xor g75 (Z[11], n_576, n_580);
  nand g76 (n_582, n_38, n_71);
  nand g77 (n_583, n_38, n_581);
  nand g78 (n_584, n_71, n_581);
  nand g79 (n_586, n_582, n_583, n_584);
  xor g80 (n_585, n_38, n_71);
  xor g81 (Z[12], n_581, n_585);
  nand g82 (n_587, n_37, n_70);
  nand g83 (n_588, n_37, n_586);
  nand g84 (n_589, n_70, n_586);
  nand g85 (n_591, n_587, n_588, n_589);
  xor g86 (n_590, n_37, n_70);
  xor g87 (Z[13], n_586, n_590);
  nand g88 (n_592, n_36, n_69);
  nand g89 (n_593, n_36, n_591);
  nand g90 (n_594, n_69, n_591);
  nand g91 (n_596, n_592, n_593, n_594);
  xor g92 (n_595, n_36, n_69);
  xor g93 (Z[14], n_591, n_595);
  nand g94 (n_597, n_35, n_68);
  nand g95 (n_598, n_35, n_596);
  nand g96 (n_599, n_68, n_596);
  nand g97 (n_601, n_597, n_598, n_599);
  xor g98 (n_600, n_35, n_68);
  xor g99 (Z[15], n_596, n_600);
  nand g552 (n_602, n_34, n_67);
  nand g553 (n_603, n_34, n_601);
  nand g554 (n_604, n_67, n_601);
  nand g555 (n_606, n_602, n_603, n_604);
  xor g556 (n_605, n_34, n_67);
  xor g557 (Z[16], n_601, n_605);
  nand g558 (n_607, n_33, n_66);
  nand g559 (n_608, n_33, n_606);
  nand g560 (n_609, n_66, n_606);
  nand g561 (n_611, n_607, n_608, n_609);
  xor g562 (n_610, n_33, n_66);
  xor g563 (Z[17], n_606, n_610);
  nand g564 (n_612, n_32, n_65);
  nand g565 (n_613, n_32, n_611);
  nand g566 (n_614, n_65, n_611);
  nand g567 (n_616, n_612, n_613, n_614);
  xor g568 (n_615, n_32, n_65);
  xor g569 (Z[18], n_611, n_615);
  nand g570 (n_617, n_31, n_64);
  nand g571 (n_618, n_31, n_616);
  nand g572 (n_619, n_64, n_616);
  nand g573 (n_621, n_617, n_618, n_619);
  xor g574 (n_620, n_31, n_64);
  xor g575 (Z[19], n_616, n_620);
  nand g576 (n_622, n_30, n_63);
  nand g577 (n_623, n_30, n_621);
  nand g578 (n_624, n_63, n_621);
  nand g579 (n_626, n_622, n_623, n_624);
  xor g580 (n_625, n_30, n_63);
  xor g581 (Z[20], n_621, n_625);
  nand g582 (n_627, n_29, n_62);
  nand g583 (n_628, n_29, n_626);
  nand g584 (n_629, n_62, n_626);
  nand g585 (n_631, n_627, n_628, n_629);
  xor g586 (n_630, n_29, n_62);
  xor g587 (Z[21], n_626, n_630);
  nand g588 (n_632, n_28, n_61);
  nand g589 (n_633, n_28, n_631);
  nand g590 (n_634, n_61, n_631);
  nand g591 (n_636, n_632, n_633, n_634);
  xor g592 (n_635, n_28, n_61);
  xor g593 (Z[22], n_631, n_635);
  nand g594 (n_637, n_27, n_60);
  nand g595 (n_638, n_27, n_636);
  nand g596 (n_639, n_60, n_636);
  nand g597 (n_641, n_637, n_638, n_639);
  xor g598 (n_640, n_27, n_60);
  xor g599 (Z[23], n_636, n_640);
  nand g600 (n_642, n_26, n_59);
  nand g601 (n_643, n_26, n_641);
  nand g602 (n_644, n_59, n_641);
  nand g603 (n_646, n_642, n_643, n_644);
  xor g604 (n_645, n_26, n_59);
  xor g605 (Z[24], n_641, n_645);
  nand g606 (n_647, n_25, n_58);
  nand g607 (n_648, n_25, n_646);
  nand g608 (n_649, n_58, n_646);
  nand g609 (n_651, n_647, n_648, n_649);
  xor g610 (n_650, n_25, n_58);
  xor g611 (Z[25], n_646, n_650);
  nand g612 (n_652, n_24, n_57);
  nand g613 (n_653, n_24, n_651);
  nand g614 (n_654, n_57, n_651);
  nand g615 (n_656, n_652, n_653, n_654);
  xor g616 (n_655, n_24, n_57);
  xor g617 (Z[26], n_651, n_655);
  nand g618 (n_657, n_23, n_56);
  nand g619 (n_658, n_23, n_656);
  nand g620 (n_659, n_56, n_656);
  nand g621 (n_661, n_657, n_658, n_659);
  xor g622 (n_660, n_23, n_56);
  xor g623 (Z[27], n_656, n_660);
  nand g624 (n_662, n_22, n_55);
  nand g625 (n_663, n_22, n_661);
  nand g626 (n_664, n_55, n_661);
  nand g627 (n_666, n_662, n_663, n_664);
  xor g628 (n_665, n_22, n_55);
  xor g629 (Z[28], n_661, n_665);
  nand g630 (n_667, n_21, n_54);
  nand g631 (n_668, n_21, n_666);
  nand g632 (n_669, n_54, n_666);
  nand g633 (n_671, n_667, n_668, n_669);
  xor g634 (n_670, n_21, n_54);
  xor g635 (Z[29], n_666, n_670);
  nand g638 (n_674, n_53, n_671);
  nand g639 (n_676, n_672, n_673, n_674);
  xor g641 (Z[30], n_671, n_675);
  nand g644 (n_679, A[15], n_676);
  nand g645 (n_681, n_677, n_678, n_679);
  xor g647 (Z[31], n_676, n_680);
  or g652 (n_122, A[4], A[6], wc);
  not gc (wc, n_253);
  or g654 (n_257, A[0], wc0);
  not gc0 (wc0, A[2]);
  xnor g655 (n_123, n_260, A[1]);
  or g656 (n_262, A[1], wc1);
  not gc1 (wc1, A[5]);
  or g657 (n_263, A[1], wc2);
  not gc2 (wc2, A[7]);
  xnor g658 (n_126, n_268, A[2]);
  or g659 (n_270, A[2], wc3);
  not gc3 (wc3, A[6]);
  or g660 (n_271, A[2], wc4);
  not gc4 (wc4, A[8]);
  xnor g661 (n_276, A[3], A[0]);
  or g662 (n_277, wc5, A[3]);
  not gc5 (wc5, A[0]);
  or g663 (n_279, A[3], wc6);
  not gc6 (wc6, A[5]);
  xnor g664 (n_134, n_284, A[4]);
  or g665 (n_286, A[4], wc7);
  not gc7 (wc7, A[8]);
  or g666 (n_287, A[4], wc8);
  not gc8 (wc8, A[10]);
  xnor g667 (n_138, n_296, A[5]);
  or g668 (n_298, A[5], wc9);
  not gc9 (wc9, A[9]);
  or g669 (n_299, A[5], wc10);
  not gc10 (wc10, A[11]);
  xnor g670 (n_143, n_308, A[6]);
  or g671 (n_310, A[6], wc11);
  not gc11 (wc11, A[10]);
  or g672 (n_311, A[6], wc12);
  not gc12 (wc12, A[12]);
  xnor g673 (n_320, A[7], A[4]);
  or g674 (n_321, wc13, A[7]);
  not gc13 (wc13, A[4]);
  or g675 (n_323, A[7], wc14);
  not gc14 (wc14, A[9]);
  xnor g676 (n_150, n_241, A[8]);
  or g677 (n_334, A[8], wc15);
  not gc15 (wc15, A[12]);
  or g678 (n_335, A[8], wc16);
  not gc16 (wc16, A[14]);
  xnor g679 (n_348, A[9], A[6]);
  or g680 (n_349, wc17, A[9]);
  not gc17 (wc17, A[6]);
  or g681 (n_351, A[9], wc18);
  not gc18 (wc18, A[11]);
  xnor g682 (n_165, A[16], A[14]);
  and g683 (n_174, A[14], wc19);
  not gc19 (wc19, A[16]);
  or g684 (n_367, wc20, A[10]);
  not gc20 (wc20, A[7]);
  xnor g685 (n_177, n_384, A[11]);
  or g686 (n_386, wc21, A[11]);
  not gc21 (wc21, A[4]);
  or g687 (n_387, wc22, A[11]);
  not gc22 (wc22, A[8]);
  xnor g688 (n_178, n_81, A[2]);
  or g691 (n_407, wc23, A[16]);
  not gc23 (wc23, A[9]);
  xnor g692 (n_408, A[12], A[5]);
  or g693 (n_409, wc24, A[12]);
  not gc24 (wc24, A[5]);
  or g694 (n_410, wc25, A[12]);
  not gc25 (wc25, A[3]);
  and g695 (n_204, wc26, A[15]);
  not gc26 (wc26, A[13]);
  or g697 (n_441, A[16], A[14]);
  or g698 (n_442, wc27, A[14]);
  not gc27 (wc27, A[7]);
  or g699 (n_443, wc28, A[16]);
  not gc28 (wc28, A[7]);
  xnor g700 (n_213, A[15], A[12]);
  and g701 (n_219, A[12], wc29);
  not gc29 (wc29, A[15]);
  or g703 (n_220, A[6], A[8], wc30);
  not gc30 (wc30, n_269);
  xnor g704 (n_227, n_225, A[8]);
  xnor g706 (n_232, n_230, A[9]);
  xnor g708 (n_496, A[16], A[12]);
  or g709 (n_497, wc31, A[16]);
  not gc31 (wc31, A[12]);
  or g710 (n_499, wc32, A[16]);
  not gc32 (wc32, A[10]);
  or g714 (n_514, wc33, n_333);
  not gc33 (wc33, n_81);
  or g715 (n_519, A[16], wc34);
  not gc34 (wc34, n_164);
  or g716 (n_677, wc35, A[16]);
  not gc35 (wc35, A[15]);
  xnor g717 (n_680, A[16], A[15]);
  xnor g718 (n_77, n_120, Z[2]);
  or g719 (n_259, A[0], wc36);
  not gc36 (wc36, n_120);
  or g720 (n_175, A[7], wc37, wc38);
  not gc38 (wc38, n_367);
  not gc37 (wc37, A[10]);
  or g721 (n_188, A[2], wc39, n_81);
  not gc39 (wc39, n_355);
  or g722 (n_197, wc40, n_174, wc41);
  not gc41 (wc41, n_406);
  not gc40 (wc40, n_407);
  xnor g723 (n_206, n_165, A[7]);
  or g724 (n_463, wc42, n_268);
  not gc42 (wc42, n_213);
  or g725 (n_233, A[8], wc43, n_225);
  not gc43 (wc43, n_482);
  or g726 (n_236, A[9], wc44, n_230);
  not gc44 (wc44, n_490);
  xnor g727 (n_56, n_148, n_241);
  or g728 (n_22, wc45, n_241, n_148);
  not gc45 (wc45, n_510);
  xor g729 (n_55, n_333, n_81);
  or g730 (n_21, wc46, n_81, wc47);
  not gc47 (wc47, n_333);
  not gc46 (wc46, n_514);
  or g731 (n_53, wc48, n_174, wc49);
  not gc49 (wc49, n_518);
  not gc48 (wc48, n_519);
  or g732 (n_430, wc50, n_81);
  not gc50 (wc50, n_196);
  or g734 (n_462, wc51, n_268);
  not gc51 (wc51, n_214);
  xnor g735 (n_24, n_47, n_239);
  or g737 (n_552, wc52, n_252);
  not gc52 (wc52, n_77);
  xnor g738 (n_555, n_252, n_77);
  or g739 (n_672, A[15], wc53);
  not gc53 (wc53, n_53);
  xnor g740 (n_675, n_53, A[15]);
  or g741 (n_208, wc54, n_196, wc55);
  not gc55 (wc55, n_81);
  not gc54 (wc54, n_430);
  xnor g742 (n_217, n_268, n_460);
  or g743 (n_23, wc56, n_239, n_47);
  not gc56 (wc56, n_506);
  or g745 (n_538, wc57, n_353);
  not gc57 (wc57, A[3]);
  or g746 (n_539, wc58, n_353);
  not gc58 (wc58, A[1]);
  xnor g747 (Z[3], n_353, n_540);
  or g748 (n_553, wc59, n_252);
  not gc59 (wc59, n_551);
  or g749 (n_673, A[15], wc60);
  not gc60 (wc60, n_671);
  or g750 (n_678, A[16], wc61);
  not gc61 (wc61, n_676);
  not g751 (Z[32], n_681);
endmodule

module mult_signed_const_608_GENERIC(A, Z);
  input [16:0] A;
  output [32:0] Z;
  wire [16:0] A;
  wire [32:0] Z;
  mult_signed_const_608_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_687_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * -1449;"
  input [16:0] A;
  output [28:0] Z;
  wire [16:0] A;
  wire [28:0] Z;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_46, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_111, n_113, n_114, n_117, n_118;
  wire n_119, n_122, n_123, n_124, n_125, n_126, n_128, n_129;
  wire n_130, n_131, n_132, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_223, n_224, n_225, n_226, n_227, n_229, n_231;
  wire n_232, n_234, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_245, n_247, n_248, n_249, n_250, n_254, n_255, n_256;
  wire n_257, n_258, n_260, n_261, n_262, n_265, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_286;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_334, n_335, n_336, n_337, n_338, n_339, n_340;
  wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_385, n_389, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_402, n_405, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_418, n_421;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_434, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_473, n_475;
  wire n_476, n_477, n_478, n_479, n_480, n_483, n_484, n_485;
  wire n_486, n_489, n_490, n_504, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567;
  wire n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575;
  wire n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591;
  wire n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599;
  wire n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615;
  wire n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_624;
  wire n_625, n_627;
  assign Z[0] = A[0];
  assign Z[27] = Z[28];
  xor g104 (n_70, A[0], n_111);
  xor g112 (n_69, n_247, n_114);
  nand g114 (n_249, n_114, n_113);
  nand g116 (n_39, n_248, n_249, n_250);
  nand g124 (n_124, A[0], A[2], n_254);
  xor g125 (n_255, n_117, n_118);
  xor g126 (n_68, n_255, n_119);
  nand g127 (n_256, n_117, n_118);
  nand g128 (n_257, n_119, n_118);
  nand g129 (n_258, n_117, n_119);
  nand g130 (n_38, n_256, n_257, n_258);
  nand g138 (n_130, n_260, n_261, n_262);
  nand g142 (n_265, n_123, n_122);
  xor g145 (n_267, n_124, n_125);
  xor g146 (n_67, n_267, n_126);
  nand g147 (n_268, n_124, n_125);
  nand g148 (n_269, n_126, n_125);
  nand g149 (n_270, n_124, n_126);
  nand g150 (n_37, n_268, n_269, n_270);
  xor g159 (n_275, n_128, n_129);
  xor g160 (n_132, n_275, n_130);
  nand g161 (n_276, n_128, n_129);
  nand g162 (n_277, n_130, n_129);
  nand g163 (n_278, n_128, n_130);
  nand g164 (n_140, n_276, n_277, n_278);
  xor g165 (n_279, n_131, n_46);
  xor g166 (n_66, n_279, n_132);
  nand g167 (n_280, n_131, n_46);
  nand g168 (n_281, n_132, n_46);
  nand g169 (n_282, n_131, n_132);
  nand g170 (n_36, n_280, n_281, n_282);
  xor g180 (n_139, A[0], n_135);
  xor g185 (n_291, n_136, n_137);
  xor g186 (n_141, n_291, n_138);
  nand g187 (n_292, n_136, n_137);
  nand g188 (n_293, n_138, n_137);
  nand g189 (n_294, n_136, n_138);
  nand g190 (n_149, n_292, n_293, n_294);
  xor g191 (n_295, n_139, n_140);
  xor g192 (n_65, n_295, n_141);
  nand g193 (n_296, n_139, n_140);
  nand g194 (n_297, n_141, n_140);
  nand g195 (n_298, n_139, n_141);
  nand g196 (n_35, n_296, n_297, n_298);
  xor g206 (n_148, n_303, n_144);
  nand g208 (n_305, n_144, n_143);
  nand g210 (n_156, n_304, n_305, n_306);
  xor g211 (n_307, n_145, n_146);
  xor g212 (n_150, n_307, n_147);
  nand g213 (n_308, n_145, n_146);
  nand g214 (n_309, n_147, n_146);
  nand g215 (n_310, n_145, n_147);
  nand g216 (n_159, n_308, n_309, n_310);
  xor g217 (n_311, n_148, n_149);
  xor g218 (n_64, n_311, n_150);
  nand g219 (n_312, n_148, n_149);
  nand g220 (n_313, n_150, n_149);
  nand g221 (n_314, n_148, n_150);
  nand g222 (n_34, n_312, n_313, n_314);
  xor g232 (n_157, n_319, n_153);
  nand g234 (n_321, n_153, n_152);
  nand g236 (n_165, n_320, n_321, n_322);
  xor g237 (n_323, n_154, n_155);
  xor g238 (n_158, n_323, n_156);
  nand g239 (n_324, n_154, n_155);
  nand g240 (n_325, n_156, n_155);
  nand g241 (n_326, n_154, n_156);
  nand g242 (n_168, n_324, n_325, n_326);
  xor g243 (n_327, n_157, n_158);
  xor g244 (n_63, n_327, n_159);
  nand g245 (n_328, n_157, n_158);
  nand g246 (n_329, n_159, n_158);
  nand g247 (n_330, n_157, n_159);
  nand g248 (n_33, n_328, n_329, n_330);
  xor g258 (n_166, n_335, n_162);
  nand g260 (n_337, n_162, n_161);
  nand g262 (n_174, n_336, n_337, n_338);
  xor g263 (n_339, n_163, n_164);
  xor g264 (n_167, n_339, n_165);
  nand g265 (n_340, n_163, n_164);
  nand g266 (n_341, n_165, n_164);
  nand g267 (n_342, n_163, n_165);
  nand g268 (n_177, n_340, n_341, n_342);
  xor g269 (n_343, n_166, n_167);
  xor g270 (n_62, n_343, n_168);
  nand g271 (n_344, n_166, n_167);
  nand g272 (n_345, n_168, n_167);
  nand g273 (n_346, n_166, n_168);
  nand g274 (n_32, n_344, n_345, n_346);
  xor g284 (n_175, n_351, n_171);
  nand g286 (n_353, n_171, n_170);
  nand g288 (n_183, n_352, n_353, n_354);
  xor g289 (n_355, n_172, n_173);
  xor g290 (n_176, n_355, n_174);
  nand g291 (n_356, n_172, n_173);
  nand g292 (n_357, n_174, n_173);
  nand g293 (n_358, n_172, n_174);
  nand g294 (n_186, n_356, n_357, n_358);
  xor g295 (n_359, n_175, n_176);
  xor g296 (n_61, n_359, n_177);
  nand g297 (n_360, n_175, n_176);
  nand g298 (n_361, n_177, n_176);
  nand g299 (n_362, n_175, n_177);
  nand g300 (n_31, n_360, n_361, n_362);
  xor g310 (n_184, n_367, n_180);
  nand g312 (n_369, n_180, n_179);
  nand g314 (n_192, n_368, n_369, n_370);
  xor g315 (n_371, n_181, n_182);
  xor g316 (n_185, n_371, n_183);
  nand g317 (n_372, n_181, n_182);
  nand g318 (n_373, n_183, n_182);
  nand g319 (n_374, n_181, n_183);
  nand g320 (n_195, n_372, n_373, n_374);
  xor g321 (n_375, n_184, n_185);
  xor g322 (n_60, n_375, n_186);
  nand g323 (n_376, n_184, n_185);
  nand g324 (n_377, n_186, n_185);
  nand g325 (n_378, n_184, n_186);
  nand g326 (n_30, n_376, n_377, n_378);
  nand g332 (n_199, n_380, n_381, n_382);
  nand g342 (n_389, n_189, n_188);
  xor g345 (n_391, n_190, n_191);
  xor g346 (n_194, n_391, n_192);
  nand g347 (n_392, n_190, n_191);
  nand g348 (n_393, n_192, n_191);
  nand g349 (n_394, n_190, n_192);
  nand g350 (n_203, n_392, n_393, n_394);
  xor g351 (n_395, n_193, n_194);
  xor g352 (n_59, n_395, n_195);
  nand g353 (n_396, n_193, n_194);
  nand g354 (n_397, n_195, n_194);
  nand g355 (n_398, n_193, n_195);
  nand g356 (n_29, n_396, n_397, n_398);
  nand g368 (n_405, n_198, n_197);
  xor g371 (n_407, n_199, n_200);
  xor g372 (n_204, n_407, n_201);
  nand g373 (n_408, n_199, n_200);
  nand g374 (n_409, n_201, n_200);
  nand g375 (n_410, n_199, n_201);
  nand g376 (n_213, n_408, n_409, n_410);
  xor g377 (n_411, n_202, n_203);
  xor g378 (n_58, n_411, n_204);
  nand g379 (n_412, n_202, n_203);
  nand g380 (n_413, n_204, n_203);
  nand g381 (n_414, n_202, n_204);
  nand g382 (n_28, n_412, n_413, n_414);
  nand g394 (n_421, n_207, n_206);
  xor g397 (n_423, n_208, n_209);
  xor g398 (n_212, n_423, n_210);
  nand g399 (n_424, n_208, n_209);
  nand g400 (n_425, n_210, n_209);
  nand g401 (n_426, n_208, n_210);
  nand g402 (n_220, n_424, n_425, n_426);
  xor g403 (n_427, n_211, n_212);
  xor g404 (n_57, n_427, n_213);
  nand g405 (n_428, n_211, n_212);
  nand g406 (n_429, n_213, n_212);
  nand g407 (n_430, n_211, n_213);
  nand g408 (n_27, n_428, n_429, n_430);
  xor g416 (n_218, n_152, n_214);
  xor g421 (n_439, n_215, n_216);
  xor g422 (n_219, n_439, n_217);
  nand g423 (n_440, n_215, n_216);
  nand g424 (n_441, n_217, n_216);
  nand g425 (n_442, n_215, n_217);
  nand g426 (n_227, n_440, n_441, n_442);
  xor g427 (n_443, n_218, n_219);
  xor g428 (n_56, n_443, n_220);
  nand g429 (n_444, n_218, n_219);
  nand g430 (n_445, n_220, n_219);
  nand g431 (n_446, n_218, n_220);
  nand g432 (n_55, n_444, n_445, n_446);
  nand g440 (n_229, A[10], A[12], n_450);
  xor g441 (n_451, n_206, n_223);
  xor g442 (n_226, n_451, n_224);
  nand g443 (n_452, n_206, n_223);
  nand g444 (n_453, n_224, n_223);
  nand g445 (n_454, n_206, n_224);
  nand g446 (n_232, n_452, n_453, n_454);
  xor g447 (n_455, n_225, n_226);
  xor g448 (n_26, n_455, n_227);
  nand g449 (n_456, n_225, n_226);
  nand g450 (n_457, n_227, n_226);
  nand g451 (n_458, n_225, n_227);
  nand g452 (n_54, n_456, n_457, n_458);
  xor g460 (n_231, n_463, n_229);
  nand g462 (n_465, n_229, n_214);
  nand g464 (n_237, n_464, n_465, n_466);
  xor g465 (n_467, n_216, n_231);
  xor g466 (n_25, n_467, n_232);
  nand g467 (n_468, n_216, n_231);
  nand g468 (n_469, n_232, n_231);
  nand g469 (n_470, n_216, n_232);
  nand g470 (n_53, n_468, n_469, n_470);
  xor g474 (n_236, A[12], n_234);
  xor g479 (n_475, n_223, n_236);
  xor g480 (n_24, n_475, n_237);
  nand g481 (n_476, n_223, n_236);
  nand g482 (n_477, n_237, n_236);
  nand g483 (n_478, n_223, n_237);
  nand g484 (n_52, n_476, n_477, n_478);
  xor g491 (n_483, n_238, n_239);
  xor g492 (n_23, n_483, n_240);
  nand g493 (n_484, n_238, n_239);
  nand g494 (n_485, n_240, n_239);
  nand g495 (n_486, n_238, n_240);
  nand g496 (n_51, n_484, n_485, n_486);
  xor g498 (n_22, n_431, n_241);
  nand g501 (n_490, A[16], n_241);
  nand g502 (n_50, n_432, n_489, n_490);
  nand g25 (n_512, n_508, n_509, n_510);
  nand g30 (n_515, n_71, n_512);
  nand g31 (n_517, n_513, n_514, n_515);
  xor g33 (Z[4], n_512, n_516);
  nand g34 (n_518, n_41, n_70);
  nand g35 (n_519, n_41, n_517);
  nand g36 (n_520, n_70, n_517);
  nand g37 (n_522, n_518, n_519, n_520);
  xor g38 (n_521, n_41, n_70);
  xor g39 (Z[5], n_517, n_521);
  nand g40 (n_523, n_40, n_69);
  nand g41 (n_524, n_40, n_522);
  nand g42 (n_525, n_69, n_522);
  nand g43 (n_527, n_523, n_524, n_525);
  xor g44 (n_526, n_40, n_69);
  xor g45 (Z[6], n_522, n_526);
  nand g46 (n_528, n_39, n_68);
  nand g47 (n_529, n_39, n_527);
  nand g48 (n_530, n_68, n_527);
  nand g49 (n_532, n_528, n_529, n_530);
  xor g50 (n_531, n_39, n_68);
  xor g51 (Z[7], n_527, n_531);
  nand g52 (n_533, n_38, n_67);
  nand g53 (n_534, n_38, n_532);
  nand g54 (n_535, n_67, n_532);
  nand g55 (n_537, n_533, n_534, n_535);
  xor g56 (n_536, n_38, n_67);
  xor g57 (Z[8], n_532, n_536);
  nand g58 (n_538, n_37, n_66);
  nand g59 (n_539, n_37, n_537);
  nand g60 (n_540, n_66, n_537);
  nand g61 (n_542, n_538, n_539, n_540);
  xor g62 (n_541, n_37, n_66);
  xor g63 (Z[9], n_537, n_541);
  nand g64 (n_543, n_36, n_65);
  nand g65 (n_544, n_36, n_542);
  nand g66 (n_545, n_65, n_542);
  nand g67 (n_547, n_543, n_544, n_545);
  xor g68 (n_546, n_36, n_65);
  xor g69 (Z[10], n_542, n_546);
  nand g70 (n_548, n_35, n_64);
  nand g71 (n_549, n_35, n_547);
  nand g72 (n_550, n_64, n_547);
  nand g73 (n_552, n_548, n_549, n_550);
  xor g74 (n_551, n_35, n_64);
  xor g75 (Z[11], n_547, n_551);
  nand g76 (n_553, n_34, n_63);
  nand g77 (n_554, n_34, n_552);
  nand g78 (n_555, n_63, n_552);
  nand g79 (n_557, n_553, n_554, n_555);
  xor g80 (n_556, n_34, n_63);
  xor g81 (Z[12], n_552, n_556);
  nand g82 (n_558, n_33, n_62);
  nand g83 (n_559, n_33, n_557);
  nand g84 (n_560, n_62, n_557);
  nand g85 (n_562, n_558, n_559, n_560);
  xor g86 (n_561, n_33, n_62);
  xor g87 (Z[13], n_557, n_561);
  nand g88 (n_563, n_32, n_61);
  nand g89 (n_564, n_32, n_562);
  nand g90 (n_565, n_61, n_562);
  nand g91 (n_567, n_563, n_564, n_565);
  xor g92 (n_566, n_32, n_61);
  xor g93 (Z[14], n_562, n_566);
  nand g94 (n_568, n_31, n_60);
  nand g95 (n_569, n_31, n_567);
  nand g96 (n_570, n_60, n_567);
  nand g520 (n_572, n_568, n_569, n_570);
  xor g521 (n_571, n_31, n_60);
  xor g522 (Z[15], n_567, n_571);
  nand g523 (n_573, n_30, n_59);
  nand g524 (n_574, n_30, n_572);
  nand g525 (n_575, n_59, n_572);
  nand g526 (n_577, n_573, n_574, n_575);
  xor g527 (n_576, n_30, n_59);
  xor g528 (Z[16], n_572, n_576);
  nand g529 (n_578, n_29, n_58);
  nand g530 (n_579, n_29, n_577);
  nand g531 (n_580, n_58, n_577);
  nand g532 (n_582, n_578, n_579, n_580);
  xor g533 (n_581, n_29, n_58);
  xor g534 (Z[17], n_577, n_581);
  nand g535 (n_583, n_28, n_57);
  nand g536 (n_584, n_28, n_582);
  nand g537 (n_585, n_57, n_582);
  nand g538 (n_587, n_583, n_584, n_585);
  xor g539 (n_586, n_28, n_57);
  xor g540 (Z[18], n_582, n_586);
  nand g541 (n_588, n_27, n_56);
  nand g542 (n_589, n_27, n_587);
  nand g543 (n_590, n_56, n_587);
  nand g544 (n_592, n_588, n_589, n_590);
  xor g545 (n_591, n_27, n_56);
  xor g546 (Z[19], n_587, n_591);
  nand g547 (n_593, n_26, n_55);
  nand g548 (n_594, n_26, n_592);
  nand g549 (n_595, n_55, n_592);
  nand g550 (n_597, n_593, n_594, n_595);
  xor g551 (n_596, n_26, n_55);
  xor g552 (Z[20], n_592, n_596);
  nand g553 (n_598, n_25, n_54);
  nand g554 (n_599, n_25, n_597);
  nand g555 (n_600, n_54, n_597);
  nand g556 (n_602, n_598, n_599, n_600);
  xor g557 (n_601, n_25, n_54);
  xor g558 (Z[21], n_597, n_601);
  nand g559 (n_603, n_24, n_53);
  nand g560 (n_604, n_24, n_602);
  nand g561 (n_605, n_53, n_602);
  nand g562 (n_607, n_603, n_604, n_605);
  xor g563 (n_606, n_24, n_53);
  xor g564 (Z[22], n_602, n_606);
  nand g565 (n_608, n_23, n_52);
  nand g566 (n_609, n_23, n_607);
  nand g567 (n_610, n_52, n_607);
  nand g568 (n_612, n_608, n_609, n_610);
  xor g569 (n_611, n_23, n_52);
  xor g570 (Z[23], n_607, n_611);
  nand g571 (n_613, n_22, n_51);
  nand g572 (n_614, n_22, n_612);
  nand g573 (n_615, n_51, n_612);
  nand g574 (n_617, n_613, n_614, n_615);
  xor g575 (n_616, n_22, n_51);
  xor g576 (Z[24], n_612, n_616);
  nand g577 (n_618, A[15], n_50);
  nand g578 (n_619, A[15], n_617);
  nand g579 (n_620, n_50, n_617);
  nand g580 (n_622, n_618, n_619, n_620);
  xor g581 (n_621, A[15], n_50);
  xor g582 (Z[25], n_617, n_621);
  nand g584 (n_624, A[16], n_622);
  nand g586 (n_627, n_480, n_624, n_625);
  xor g588 (Z[26], n_622, n_479);
  xor g597 (n_71, A[4], A[1]);
  nor g598 (n_41, A[4], A[1]);
  xor g599 (n_111, A[5], A[2]);
  nor g600 (n_114, A[5], A[2]);
  xor g601 (n_113, A[6], A[3]);
  nor g602 (n_118, A[6], A[3]);
  xor g603 (n_117, A[7], A[4]);
  nor g604 (n_123, A[7], A[4]);
  or g605 (n_254, A[2], A[0]);
  xor g606 (n_122, A[8], A[5]);
  nor g607 (n_129, A[8], A[5]);
  xor g608 (Z[1], A[1], A[0]);
  or g609 (n_260, A[1], A[0]);
  or g610 (n_261, A[3], A[0]);
  or g611 (n_262, A[3], A[1]);
  xor g612 (n_128, A[9], A[6]);
  nor g613 (n_135, A[9], A[6]);
  xor g614 (n_271, A[2], A[1]);
  or g615 (n_272, A[2], A[1]);
  or g617 (n_274, A[4], A[2]);
  xor g618 (n_136, A[10], A[7]);
  nor g619 (n_144, A[10], A[7]);
  xor g620 (n_283, A[3], A[2]);
  or g621 (n_284, A[3], A[2]);
  or g623 (n_286, A[5], A[3]);
  xor g624 (n_143, A[11], A[8]);
  nor g625 (n_153, A[11], A[8]);
  xor g626 (n_299, A[4], A[3]);
  or g627 (n_300, A[4], A[3]);
  or g629 (n_302, A[6], A[4]);
  xor g630 (n_152, A[12], A[9]);
  nor g631 (n_162, A[12], A[9]);
  xor g632 (n_315, A[5], A[4]);
  or g633 (n_316, A[5], A[4]);
  or g635 (n_318, A[7], A[5]);
  xor g636 (n_161, A[13], A[10]);
  nor g637 (n_171, A[13], A[10]);
  xor g638 (n_331, A[6], A[5]);
  or g639 (n_332, A[6], A[5]);
  or g641 (n_334, A[8], A[6]);
  xor g642 (n_170, A[14], A[11]);
  nor g643 (n_180, A[14], A[11]);
  xor g644 (n_347, A[7], A[6]);
  or g645 (n_348, A[7], A[6]);
  or g647 (n_350, A[9], A[7]);
  xor g648 (n_179, A[15], A[12]);
  nor g649 (n_188, A[15], A[12]);
  xor g650 (n_363, A[8], A[7]);
  or g651 (n_364, A[8], A[7]);
  or g653 (n_366, A[10], A[8]);
  xnor g654 (n_379, A[16], A[13]);
  or g655 (n_380, A[13], wc);
  not gc (wc, A[16]);
  or g656 (n_381, A[13], A[9]);
  or g657 (n_382, A[9], wc0);
  not gc0 (wc0, A[16]);
  or g659 (n_385, A[11], A[6]);
  xor g660 (n_197, A[14], A[12]);
  nor g661 (n_207, A[14], A[12]);
  xor g662 (n_399, A[9], A[7]);
  or g663 (n_402, A[10], A[9]);
  xor g664 (n_206, A[15], A[13]);
  nor g665 (n_214, A[15], A[13]);
  xor g666 (n_415, A[10], A[8]);
  or g667 (n_418, A[11], A[10]);
  xnor g668 (n_431, A[16], A[14]);
  or g669 (n_432, A[14], wc1);
  not gc1 (wc1, A[16]);
  or g671 (n_434, A[11], wc2);
  not gc2 (wc2, A[16]);
  or g673 (n_450, A[12], A[10]);
  xor g674 (n_234, A[15], A[14]);
  nor g675 (n_238, A[15], A[14]);
  xnor g676 (n_479, A[16], A[15]);
  or g677 (n_480, A[15], wc3);
  not gc3 (wc3, A[16]);
  or g679 (n_245, A[0], wc4);
  not gc4 (wc4, n_111);
  xnor g681 (n_247, n_113, A[1]);
  or g682 (n_248, A[1], wc5);
  not gc5 (wc5, n_113);
  or g683 (n_250, A[1], wc6);
  not gc6 (wc6, n_114);
  xnor g684 (n_119, A[2], A[0]);
  xnor g685 (n_125, Z[1], A[3]);
  xnor g687 (n_131, n_271, A[4]);
  or g688 (n_137, wc7, wc8, n_41);
  not gc8 (wc8, n_272);
  not gc7 (wc7, n_274);
  xnor g689 (n_138, n_283, A[5]);
  or g690 (n_145, wc9, wc10, n_114);
  not gc10 (wc10, n_284);
  not gc9 (wc9, n_286);
  or g691 (n_290, A[0], wc11);
  not gc11 (wc11, n_135);
  xnor g692 (n_146, n_299, A[6]);
  or g693 (n_154, wc12, wc13, n_118);
  not gc13 (wc13, n_300);
  not gc12 (wc12, n_302);
  xnor g694 (n_303, n_143, A[1]);
  or g695 (n_304, A[1], wc14);
  not gc14 (wc14, n_143);
  or g696 (n_306, A[1], wc15);
  not gc15 (wc15, n_144);
  xnor g697 (n_155, n_315, A[7]);
  or g698 (n_163, wc16, wc17, n_123);
  not gc17 (wc17, n_316);
  not gc16 (wc16, n_318);
  xnor g699 (n_319, n_152, A[2]);
  or g700 (n_320, A[2], wc18);
  not gc18 (wc18, n_152);
  or g701 (n_322, A[2], wc19);
  not gc19 (wc19, n_153);
  xnor g702 (n_164, n_331, A[8]);
  or g703 (n_172, wc20, wc21, n_129);
  not gc21 (wc21, n_332);
  not gc20 (wc20, n_334);
  xnor g704 (n_335, n_161, A[3]);
  or g705 (n_336, A[3], wc22);
  not gc22 (wc22, n_161);
  or g706 (n_338, A[3], wc23);
  not gc23 (wc23, n_162);
  xnor g707 (n_173, n_347, A[9]);
  or g708 (n_181, wc24, wc25, n_135);
  not gc25 (wc25, n_348);
  not gc24 (wc24, n_350);
  xnor g709 (n_351, n_170, A[4]);
  or g710 (n_352, A[4], wc26);
  not gc26 (wc26, n_170);
  or g711 (n_354, A[4], wc27);
  not gc27 (wc27, n_171);
  xnor g712 (n_182, n_363, A[10]);
  or g713 (n_189, wc28, wc29, n_144);
  not gc29 (wc29, n_364);
  not gc28 (wc28, n_366);
  xnor g714 (n_367, n_179, A[5]);
  or g715 (n_368, A[5], wc30);
  not gc30 (wc30, n_179);
  or g716 (n_370, A[5], wc31);
  not gc31 (wc31, n_180);
  xnor g717 (n_191, n_379, A[9]);
  xnor g718 (n_190, n_143, A[6]);
  or g719 (n_198, wc32, wc33, n_153);
  not gc33 (wc33, n_334);
  not gc32 (wc32, n_385);
  xnor g721 (n_200, n_399, A[10]);
  or g722 (n_208, wc34, wc35, n_144);
  not gc35 (wc35, n_350);
  not gc34 (wc34, n_402);
  xnor g724 (n_209, n_415, A[11]);
  or g725 (n_215, wc36, wc37, n_153);
  not gc37 (wc37, n_366);
  not gc36 (wc36, n_418);
  xnor g728 (n_216, n_431, A[11]);
  or g729 (n_223, wc38, wc39, n_180);
  not gc39 (wc39, n_432);
  not gc38 (wc38, n_434);
  or g730 (n_437, A[12], wc40);
  not gc40 (wc40, n_214);
  or g731 (n_438, A[9], wc41);
  not gc41 (wc41, n_214);
  xnor g732 (n_224, A[12], A[10]);
  xnor g733 (n_463, n_214, A[13]);
  or g734 (n_464, A[13], wc42);
  not gc42 (wc42, n_214);
  or g735 (n_473, A[12], wc43);
  not gc43 (wc43, n_234);
  xnor g737 (n_239, n_479, A[13]);
  or g738 (n_241, wc44, n_214, wc45);
  not gc45 (wc45, n_380);
  not gc44 (wc44, n_480);
  or g739 (n_508, A[0], wc46);
  not gc46 (wc46, A[3]);
  xnor g740 (n_511, A[3], A[0]);
  or g741 (n_513, A[3], wc47);
  not gc47 (wc47, n_71);
  xnor g742 (n_516, n_71, A[3]);
  or g743 (n_40, wc48, wc49, n_111);
  not gc49 (wc49, n_245);
  not gc48 (wc48, A[0]);
  xnor g744 (n_126, n_123, n_122);
  or g745 (n_46, n_122, n_123, wc50);
  not gc50 (wc50, n_265);
  or g746 (n_147, wc51, wc52, n_135);
  not gc52 (wc52, n_290);
  not gc51 (wc51, A[0]);
  xnor g747 (n_193, n_188, n_189);
  xnor g749 (n_201, n_197, n_198);
  xnor g751 (n_210, n_207, n_206);
  or g752 (n_217, n_206, n_207, wc53);
  not gc53 (wc53, n_421);
  or g753 (n_225, wc54, wc55, n_162);
  not gc55 (wc55, n_437);
  not gc54 (wc54, n_438);
  or g754 (n_466, A[13], wc56);
  not gc56 (wc56, n_229);
  or g755 (n_240, wc57, wc58, n_234);
  not gc58 (wc58, n_473);
  not gc57 (wc57, A[12]);
  or g756 (n_489, A[14], wc59);
  not gc59 (wc59, n_241);
  or g757 (n_202, n_189, n_188, wc60);
  not gc60 (wc60, n_389);
  or g758 (n_211, n_198, n_197, wc61);
  not gc61 (wc61, n_405);
  or g760 (n_504, n_260, A[2]);
  xor g761 (Z[2], n_260, A[2]);
  or g763 (n_509, n_504, A[0]);
  or g764 (n_510, wc62, n_504);
  not gc62 (wc62, A[3]);
  xnor g765 (Z[3], n_511, n_504);
  or g766 (n_514, A[3], wc63);
  not gc63 (wc63, n_512);
  or g767 (n_625, A[15], wc64);
  not gc64 (wc64, n_622);
  not g768 (Z[28], n_627);
endmodule

module mult_signed_const_687_GENERIC(A, Z);
  input [16:0] A;
  output [28:0] Z;
  wire [16:0] A;
  wire [28:0] Z;
  mult_signed_const_687_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_751_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 1899;"
  input [16:0] A;
  output [27:0] Z;
  wire [16:0] A;
  wire [27:0] Z;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_41, n_42, n_43, n_45, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_72, n_105, n_107, n_108;
  wire n_111, n_112, n_113, n_115, n_116, n_117, n_118, n_120;
  wire n_121, n_122, n_123, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_132, n_133, n_134, n_135, n_136, n_137, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_176, n_177;
  wire n_179, n_180, n_181, n_183, n_184, n_185, n_186, n_187;
  wire n_191, n_192, n_193, n_194, n_196, n_198, n_199, n_200;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_230, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_273, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_351, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_406, n_408, n_409, n_410, n_411;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_422;
  wire n_424, n_425, n_426, n_427, n_435, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_559, n_560, n_561, n_562, n_564;
  assign Z[0] = A[0];
  xor g83 (n_70, A[3], A[0]);
  and g84 (n_41, A[3], A[0]);
  xor g85 (n_204, A[4], A[3]);
  xor g86 (n_69, n_204, A[1]);
  nand g87 (n_205, A[4], A[3]);
  nand g88 (n_206, A[1], A[3]);
  nand g89 (n_207, A[4], A[1]);
  nand g90 (n_105, n_205, n_206, n_207);
  xor g91 (n_208, A[5], A[4]);
  nand g93 (n_209, A[5], A[4]);
  xor g98 (n_68, n_212, n_105);
  nand g100 (n_214, n_105, A[2]);
  nand g102 (n_39, n_213, n_214, n_215);
  xor g103 (n_216, A[6], A[5]);
  nand g105 (n_217, A[6], A[5]);
  nand g108 (n_111, n_217, n_218, n_219);
  xor g109 (n_220, A[3], n_107);
  xor g110 (n_67, n_220, n_108);
  nand g111 (n_221, A[3], n_107);
  nand g112 (n_222, n_108, n_107);
  nand g113 (n_223, A[3], n_108);
  nand g114 (n_38, n_221, n_222, n_223);
  xor g115 (n_224, A[7], A[6]);
  nand g117 (n_225, A[7], A[6]);
  nand g120 (n_116, n_225, n_226, n_227);
  xor g122 (n_112, A[0], A[4]);
  xor g127 (n_232, n_111, n_112);
  xor g128 (n_66, n_232, n_113);
  nand g129 (n_233, n_111, n_112);
  nand g130 (n_234, n_113, n_112);
  nand g131 (n_235, n_111, n_113);
  nand g132 (n_37, n_233, n_234, n_235);
  xor g133 (n_236, A[8], A[7]);
  nand g135 (n_237, A[8], A[7]);
  nand g138 (n_120, n_237, n_238, n_239);
  xor g140 (n_118, n_240, n_115);
  nand g142 (n_242, n_115, A[5]);
  nand g144 (n_123, n_218, n_242, n_243);
  xor g145 (n_244, n_116, n_117);
  xor g146 (n_65, n_244, n_118);
  nand g147 (n_245, n_116, n_117);
  nand g148 (n_246, n_118, n_117);
  nand g149 (n_247, n_116, n_118);
  nand g150 (n_36, n_245, n_246, n_247);
  xor g151 (n_248, A[9], A[8]);
  nand g153 (n_249, A[9], A[8]);
  nand g156 (n_125, n_249, n_250, n_251);
  xor g158 (n_122, n_252, n_120);
  nand g160 (n_254, n_120, A[6]);
  nand g162 (n_43, n_226, n_254, n_255);
  xor g163 (n_256, n_121, n_122);
  xor g164 (n_64, n_256, n_123);
  nand g165 (n_257, n_121, n_122);
  nand g166 (n_258, n_123, n_122);
  nand g167 (n_259, n_121, n_123);
  nand g168 (n_35, n_257, n_258, n_259);
  xor g169 (n_260, A[10], A[9]);
  nand g171 (n_261, A[10], A[9]);
  nand g174 (n_127, n_261, n_262, n_263);
  xor g176 (n_42, n_264, n_125);
  nand g178 (n_266, n_125, A[7]);
  nand g180 (n_130, n_238, n_266, n_267);
  xor g181 (n_268, n_126, n_42);
  xor g182 (n_63, n_268, n_43);
  nand g183 (n_269, n_126, n_42);
  nand g184 (n_270, n_43, n_42);
  nand g185 (n_271, n_126, n_43);
  nand g186 (n_34, n_269, n_270, n_271);
  xor g187 (n_45, A[11], A[10]);
  and g188 (n_132, A[11], A[10]);
  xor g190 (n_128, n_272, A[8]);
  nand g194 (n_133, n_273, n_250, n_275);
  xor g195 (n_276, A[0], n_45);
  xor g196 (n_129, n_276, n_127);
  nand g197 (n_277, A[0], n_45);
  nand g198 (n_278, n_127, n_45);
  nand g199 (n_279, A[0], n_127);
  nand g200 (n_136, n_277, n_278, n_279);
  xor g201 (n_280, n_128, n_129);
  xor g202 (n_62, n_280, n_130);
  nand g203 (n_281, n_128, n_129);
  nand g204 (n_282, n_130, n_129);
  nand g205 (n_283, n_128, n_130);
  nand g206 (n_33, n_281, n_282, n_283);
  xor g207 (n_284, A[12], A[11]);
  nand g209 (n_285, A[12], A[11]);
  nand g212 (n_140, n_285, n_286, n_287);
  xor g214 (n_135, n_288, A[1]);
  nand g216 (n_290, A[1], A[9]);
  nand g218 (n_139, n_262, n_290, n_291);
  xor g219 (n_292, n_132, n_133);
  xor g220 (n_137, n_292, n_134);
  nand g221 (n_293, n_132, n_133);
  nand g222 (n_294, n_134, n_133);
  nand g223 (n_295, n_132, n_134);
  nand g224 (n_144, n_293, n_294, n_295);
  xor g225 (n_296, n_135, n_136);
  xor g226 (n_61, n_296, n_137);
  nand g227 (n_297, n_135, n_136);
  nand g228 (n_298, n_137, n_136);
  nand g229 (n_299, n_135, n_137);
  nand g230 (n_32, n_297, n_298, n_299);
  xor g231 (n_300, A[13], A[12]);
  nand g233 (n_301, A[13], A[12]);
  nand g236 (n_147, n_301, n_302, n_303);
  xor g238 (n_142, n_304, A[2]);
  nand g240 (n_306, A[2], A[10]);
  nand g242 (n_146, n_305, n_306, n_307);
  xor g243 (n_308, n_139, n_140);
  xor g244 (n_143, n_308, n_141);
  nand g245 (n_309, n_139, n_140);
  nand g246 (n_310, n_141, n_140);
  nand g247 (n_311, n_139, n_141);
  nand g248 (n_151, n_309, n_310, n_311);
  xor g249 (n_312, n_142, n_143);
  xor g250 (n_60, n_312, n_144);
  nand g251 (n_313, n_142, n_143);
  nand g252 (n_314, n_144, n_143);
  nand g253 (n_315, n_142, n_144);
  nand g254 (n_31, n_313, n_314, n_315);
  xor g255 (n_316, A[14], A[13]);
  nand g257 (n_317, A[14], A[13]);
  nand g260 (n_152, n_317, n_318, n_319);
  xor g262 (n_149, n_320, A[3]);
  nand g264 (n_322, A[3], A[11]);
  nand g266 (n_72, n_286, n_322, n_323);
  xor g267 (n_324, n_146, n_147);
  xor g268 (n_150, n_324, n_148);
  nand g269 (n_325, n_146, n_147);
  nand g270 (n_326, n_148, n_147);
  nand g271 (n_327, n_146, n_148);
  nand g272 (n_156, n_325, n_326, n_327);
  xor g273 (n_328, n_149, n_150);
  xor g274 (n_59, n_328, n_151);
  nand g275 (n_329, n_149, n_150);
  nand g276 (n_330, n_151, n_150);
  nand g277 (n_331, n_149, n_151);
  nand g278 (n_30, n_329, n_330, n_331);
  xor g279 (n_332, A[15], A[14]);
  nand g281 (n_333, A[15], A[14]);
  nand g284 (n_160, n_333, n_334, n_335);
  xor g286 (n_154, n_336, A[4]);
  nand g288 (n_338, A[4], A[12]);
  nand g290 (n_161, n_302, n_338, n_339);
  xor g291 (n_340, n_72, n_152);
  xor g292 (n_155, n_340, n_153);
  nand g293 (n_341, n_72, n_152);
  nand g294 (n_342, n_153, n_152);
  nand g295 (n_343, n_72, n_153);
  nand g296 (n_165, n_341, n_342, n_343);
  xor g297 (n_344, n_154, n_155);
  xor g298 (n_58, n_344, n_156);
  nand g299 (n_345, n_154, n_155);
  nand g300 (n_346, n_156, n_155);
  nand g301 (n_347, n_154, n_156);
  nand g302 (n_29, n_345, n_346, n_347);
  xor g306 (n_162, n_348, A[13]);
  nand g310 (n_168, n_349, n_318, n_351);
  nand g315 (n_355, A[5], n_159);
  xor g317 (n_356, n_160, n_161);
  xor g318 (n_164, n_356, n_162);
  nand g319 (n_357, n_160, n_161);
  nand g320 (n_358, n_162, n_161);
  nand g321 (n_359, n_160, n_162);
  nand g322 (n_172, n_357, n_358, n_359);
  xor g323 (n_360, n_163, n_164);
  xor g324 (n_57, n_360, n_165);
  nand g325 (n_361, n_163, n_164);
  nand g326 (n_362, n_165, n_164);
  nand g327 (n_363, n_163, n_165);
  nand g328 (n_28, n_361, n_362, n_363);
  nand g334 (n_177, n_365, n_334, n_367);
  xor g336 (n_171, n_368, n_167);
  nand g339 (n_371, A[6], n_167);
  nand g340 (n_179, n_369, n_370, n_371);
  xor g341 (n_372, n_168, n_169);
  xor g342 (n_173, n_372, n_170);
  nand g343 (n_373, n_168, n_169);
  nand g344 (n_374, n_170, n_169);
  nand g345 (n_375, n_168, n_170);
  nand g346 (n_181, n_373, n_374, n_375);
  xor g347 (n_376, n_171, n_172);
  xor g348 (n_56, n_376, n_173);
  nand g349 (n_377, n_171, n_172);
  nand g350 (n_378, n_173, n_172);
  nand g351 (n_379, n_171, n_173);
  nand g352 (n_27, n_377, n_378, n_379);
  xor g361 (n_384, n_176, n_177);
  nand g363 (n_385, n_176, n_177);
  nand g366 (n_187, n_385, n_386, n_387);
  xor g367 (n_388, n_179, n_180);
  xor g368 (n_55, n_388, n_181);
  nand g369 (n_389, n_179, n_180);
  nand g370 (n_390, n_181, n_180);
  nand g371 (n_391, n_179, n_181);
  nand g372 (n_54, n_389, n_390, n_391);
  nand g378 (n_191, n_393, n_394, n_395);
  xor g380 (n_186, n_396, n_184);
  nand g382 (n_398, n_184, n_183);
  nand g384 (n_193, n_397, n_398, n_399);
  xor g385 (n_400, n_185, n_186);
  xor g386 (n_26, n_400, n_187);
  nand g387 (n_401, n_185, n_186);
  nand g388 (n_402, n_187, n_186);
  nand g389 (n_403, n_185, n_187);
  nand g390 (n_53, n_401, n_402, n_403);
  xor g399 (n_408, n_191, n_192);
  xor g400 (n_25, n_408, n_193);
  nand g401 (n_409, n_191, n_192);
  nand g402 (n_410, n_193, n_192);
  nand g403 (n_411, n_191, n_193);
  nand g404 (n_52, n_409, n_410, n_411);
  nand g409 (n_415, A[16], A[10]);
  nand g410 (n_199, n_413, n_414, n_415);
  xor g412 (n_24, n_416, n_196);
  nand g415 (n_419, n_194, n_196);
  nand g416 (n_51, n_417, n_418, n_419);
  nand g422 (n_422, n_199, n_198);
  xor g425 (n_424, A[16], A[12]);
  xor g426 (n_22, n_424, n_200);
  nand g427 (n_425, A[16], A[12]);
  nand g428 (n_426, n_200, A[12]);
  nand g429 (n_427, A[16], n_200);
  nand g430 (n_49, n_425, n_426, n_427);
  nand g445 (n_435, A[1], A[0]);
  xor g449 (Z[1], A[1], A[0]);
  nand g451 (n_440, A[2], A[1]);
  nand g19 (n_444, n_440, n_441, n_442);
  xor g20 (n_443, A[2], A[1]);
  nand g22 (n_445, A[2], n_70);
  nand g23 (n_446, A[2], n_444);
  nand g24 (n_447, n_70, n_444);
  nand g25 (n_449, n_445, n_446, n_447);
  xor g26 (n_448, A[2], n_70);
  xor g27 (Z[3], n_444, n_448);
  nand g28 (n_450, n_41, n_69);
  nand g29 (n_451, n_41, n_449);
  nand g30 (n_452, n_69, n_449);
  nand g31 (n_454, n_450, n_451, n_452);
  xor g32 (n_453, n_41, n_69);
  xor g33 (Z[4], n_449, n_453);
  nand g36 (n_457, n_68, n_454);
  nand g37 (n_459, n_455, n_456, n_457);
  xor g39 (Z[5], n_454, n_458);
  nand g40 (n_460, n_39, n_67);
  nand g41 (n_461, n_39, n_459);
  nand g42 (n_462, n_67, n_459);
  nand g43 (n_464, n_460, n_461, n_462);
  xor g44 (n_463, n_39, n_67);
  xor g45 (Z[6], n_459, n_463);
  nand g46 (n_465, n_38, n_66);
  nand g47 (n_466, n_38, n_464);
  nand g48 (n_467, n_66, n_464);
  nand g49 (n_469, n_465, n_466, n_467);
  xor g50 (n_468, n_38, n_66);
  xor g51 (Z[7], n_464, n_468);
  nand g52 (n_470, n_37, n_65);
  nand g53 (n_471, n_37, n_469);
  nand g54 (n_472, n_65, n_469);
  nand g55 (n_474, n_470, n_471, n_472);
  xor g56 (n_473, n_37, n_65);
  xor g57 (Z[8], n_469, n_473);
  nand g58 (n_475, n_36, n_64);
  nand g59 (n_476, n_36, n_474);
  nand g60 (n_477, n_64, n_474);
  nand g61 (n_479, n_475, n_476, n_477);
  xor g62 (n_478, n_36, n_64);
  xor g63 (Z[9], n_474, n_478);
  nand g64 (n_480, n_35, n_63);
  nand g65 (n_481, n_35, n_479);
  nand g66 (n_482, n_63, n_479);
  nand g67 (n_484, n_480, n_481, n_482);
  xor g68 (n_483, n_35, n_63);
  xor g69 (Z[10], n_479, n_483);
  nand g70 (n_485, n_34, n_62);
  nand g71 (n_486, n_34, n_484);
  nand g72 (n_487, n_62, n_484);
  nand g73 (n_489, n_485, n_486, n_487);
  xor g74 (n_488, n_34, n_62);
  xor g75 (Z[11], n_484, n_488);
  nand g76 (n_490, n_33, n_61);
  nand g77 (n_491, n_33, n_489);
  nand g78 (n_492, n_61, n_489);
  nand g79 (n_494, n_490, n_491, n_492);
  xor g80 (n_493, n_33, n_61);
  xor g81 (Z[12], n_489, n_493);
  nand g82 (n_495, n_32, n_60);
  nand g453 (n_496, n_32, n_494);
  nand g454 (n_497, n_60, n_494);
  nand g455 (n_499, n_495, n_496, n_497);
  xor g456 (n_498, n_32, n_60);
  xor g457 (Z[13], n_494, n_498);
  nand g458 (n_500, n_31, n_59);
  nand g459 (n_501, n_31, n_499);
  nand g460 (n_502, n_59, n_499);
  nand g461 (n_504, n_500, n_501, n_502);
  xor g462 (n_503, n_31, n_59);
  xor g463 (Z[14], n_499, n_503);
  nand g464 (n_505, n_30, n_58);
  nand g465 (n_506, n_30, n_504);
  nand g466 (n_507, n_58, n_504);
  nand g467 (n_509, n_505, n_506, n_507);
  xor g468 (n_508, n_30, n_58);
  xor g469 (Z[15], n_504, n_508);
  nand g470 (n_510, n_29, n_57);
  nand g471 (n_511, n_29, n_509);
  nand g472 (n_512, n_57, n_509);
  nand g473 (n_514, n_510, n_511, n_512);
  xor g474 (n_513, n_29, n_57);
  xor g475 (Z[16], n_509, n_513);
  nand g476 (n_515, n_28, n_56);
  nand g477 (n_516, n_28, n_514);
  nand g478 (n_517, n_56, n_514);
  nand g479 (n_519, n_515, n_516, n_517);
  xor g480 (n_518, n_28, n_56);
  xor g481 (Z[17], n_514, n_518);
  nand g482 (n_520, n_27, n_55);
  nand g483 (n_521, n_27, n_519);
  nand g484 (n_522, n_55, n_519);
  nand g485 (n_524, n_520, n_521, n_522);
  xor g486 (n_523, n_27, n_55);
  xor g487 (Z[18], n_519, n_523);
  nand g488 (n_525, n_26, n_54);
  nand g489 (n_526, n_26, n_524);
  nand g490 (n_527, n_54, n_524);
  nand g491 (n_529, n_525, n_526, n_527);
  xor g492 (n_528, n_26, n_54);
  xor g493 (Z[19], n_524, n_528);
  nand g494 (n_530, n_25, n_53);
  nand g495 (n_531, n_25, n_529);
  nand g496 (n_532, n_53, n_529);
  nand g497 (n_534, n_530, n_531, n_532);
  xor g498 (n_533, n_25, n_53);
  xor g499 (Z[20], n_529, n_533);
  nand g500 (n_535, n_24, n_52);
  nand g501 (n_536, n_24, n_534);
  nand g502 (n_537, n_52, n_534);
  nand g503 (n_539, n_535, n_536, n_537);
  xor g504 (n_538, n_24, n_52);
  xor g505 (Z[21], n_534, n_538);
  nand g506 (n_540, n_23, n_51);
  nand g507 (n_541, n_23, n_539);
  nand g508 (n_542, n_51, n_539);
  nand g509 (n_544, n_540, n_541, n_542);
  xor g510 (n_543, n_23, n_51);
  xor g511 (Z[22], n_539, n_543);
  nand g512 (n_545, n_22, n_50);
  nand g513 (n_546, n_22, n_544);
  nand g514 (n_547, n_50, n_544);
  nand g515 (n_549, n_545, n_546, n_547);
  xor g516 (n_548, n_22, n_50);
  xor g517 (Z[23], n_544, n_548);
  nand g520 (n_552, n_49, n_549);
  nand g521 (n_554, n_550, n_551, n_552);
  xor g523 (Z[24], n_549, n_553);
  nand g525 (n_556, A[13], n_554);
  nand g527 (n_559, n_555, n_556, n_557);
  nand g531 (n_561, A[14], n_559);
  nand g533 (n_564, n_560, n_561, n_562);
  xor g537 (Z[27], n_564, n_159);
  or g539 (n_107, A[4], A[5], wc);
  not gc (wc, n_209);
  xnor g540 (n_212, A[2], A[0]);
  or g541 (n_213, A[0], wc0);
  not gc0 (wc0, A[2]);
  xnor g542 (n_108, n_216, A[1]);
  or g543 (n_218, A[1], wc1);
  not gc1 (wc1, A[5]);
  or g544 (n_219, A[1], wc2);
  not gc2 (wc2, A[6]);
  xnor g545 (n_113, n_224, A[2]);
  or g546 (n_226, A[2], wc3);
  not gc3 (wc3, A[6]);
  or g547 (n_227, A[2], wc4);
  not gc4 (wc4, A[7]);
  or g548 (n_230, A[0], wc5);
  not gc5 (wc5, A[4]);
  xnor g549 (n_117, n_236, A[3]);
  or g550 (n_238, A[3], wc6);
  not gc6 (wc6, A[7]);
  or g551 (n_239, A[3], wc7);
  not gc7 (wc7, A[8]);
  xnor g552 (n_240, A[5], A[1]);
  xnor g553 (n_121, n_248, A[4]);
  or g554 (n_250, A[4], wc8);
  not gc8 (wc8, A[8]);
  or g555 (n_251, A[4], wc9);
  not gc9 (wc9, A[9]);
  xnor g556 (n_252, A[6], A[2]);
  xnor g557 (n_126, n_260, A[5]);
  or g558 (n_262, A[5], wc10);
  not gc10 (wc10, A[9]);
  or g559 (n_263, A[5], wc11);
  not gc11 (wc11, A[10]);
  xnor g560 (n_264, A[7], A[3]);
  xor g561 (n_272, A[6], A[4]);
  or g562 (n_273, A[6], A[4]);
  or g563 (n_275, A[6], wc12);
  not gc12 (wc12, A[8]);
  xnor g564 (n_134, n_284, A[7]);
  or g565 (n_286, A[7], wc13);
  not gc13 (wc13, A[11]);
  or g566 (n_287, A[7], wc14);
  not gc14 (wc14, A[12]);
  xnor g567 (n_288, A[9], A[5]);
  or g568 (n_291, wc15, A[5]);
  not gc15 (wc15, A[1]);
  xnor g569 (n_141, n_300, A[8]);
  or g570 (n_302, A[8], wc16);
  not gc16 (wc16, A[12]);
  or g571 (n_303, A[8], wc17);
  not gc17 (wc17, A[13]);
  xnor g572 (n_304, A[10], A[6]);
  or g573 (n_305, A[6], wc18);
  not gc18 (wc18, A[10]);
  or g574 (n_307, wc19, A[6]);
  not gc19 (wc19, A[2]);
  xnor g575 (n_148, n_316, A[9]);
  or g576 (n_318, A[9], wc20);
  not gc20 (wc20, A[13]);
  or g577 (n_319, A[9], wc21);
  not gc21 (wc21, A[14]);
  xnor g578 (n_320, A[11], A[7]);
  or g579 (n_323, wc22, A[7]);
  not gc22 (wc22, A[3]);
  xnor g580 (n_153, n_332, A[10]);
  or g581 (n_334, A[10], wc23);
  not gc23 (wc23, A[14]);
  or g582 (n_335, A[10], wc24);
  not gc24 (wc24, A[15]);
  xnor g583 (n_336, A[12], A[8]);
  or g584 (n_339, wc25, A[8]);
  not gc25 (wc25, A[4]);
  xnor g585 (n_159, A[16], A[15]);
  and g586 (n_167, A[15], wc26);
  not gc26 (wc26, A[16]);
  xor g587 (n_348, A[11], A[9]);
  or g588 (n_349, A[11], A[9]);
  or g589 (n_351, A[11], wc27);
  not gc27 (wc27, A[13]);
  xnor g590 (n_364, A[16], A[14]);
  or g591 (n_365, wc28, A[16]);
  not gc28 (wc28, A[14]);
  or g592 (n_367, A[16], A[10]);
  xnor g593 (n_368, A[12], A[6]);
  or g594 (n_369, wc29, A[12]);
  not gc29 (wc29, A[6]);
  xnor g595 (n_176, A[15], A[13]);
  and g596 (n_183, wc30, A[15]);
  not gc30 (wc30, A[13]);
  or g598 (n_383, wc31, A[11]);
  not gc31 (wc31, A[7]);
  or g600 (n_393, A[16], A[14]);
  or g601 (n_394, wc32, A[14]);
  not gc32 (wc32, A[8]);
  or g602 (n_395, wc33, A[16]);
  not gc33 (wc33, A[8]);
  nor g604 (n_194, A[15], A[13]);
  or g605 (n_413, A[14], wc34);
  not gc34 (wc34, A[16]);
  or g606 (n_414, wc35, A[14]);
  not gc35 (wc35, A[10]);
  xnor g607 (n_198, A[15], A[11]);
  and g608 (n_200, A[11], wc36);
  not gc36 (wc36, A[15]);
  or g609 (n_555, wc37, A[14]);
  not gc37 (wc37, A[13]);
  or g611 (n_560, wc38, A[15]);
  not gc38 (wc38, A[14]);
  or g613 (n_215, A[0], wc39);
  not gc39 (wc39, n_105);
  or g614 (n_115, wc40, A[4], wc41);
  not gc41 (wc41, n_230);
  not gc40 (wc40, A[0]);
  xnor g615 (n_163, n_159, A[5]);
  xnor g617 (n_169, n_364, A[10]);
  or g618 (n_370, A[12], wc42);
  not gc42 (wc42, n_167);
  or g619 (n_184, A[7], wc43, wc44);
  not gc44 (wc44, n_383);
  not gc43 (wc43, A[11]);
  or g620 (n_387, wc45, n_320);
  not gc45 (wc45, n_176);
  xnor g621 (n_185, n_364, A[8]);
  xnor g622 (n_396, n_183, A[12]);
  or g623 (n_397, A[12], wc46);
  not gc46 (wc46, n_183);
  xor g624 (n_192, n_176, A[9]);
  or g625 (n_406, wc47, n_176);
  not gc47 (wc47, A[9]);
  or g628 (n_243, A[1], wc48);
  not gc48 (wc48, n_115);
  or g629 (n_255, A[2], wc49);
  not gc49 (wc49, n_120);
  or g630 (n_267, A[3], wc50);
  not gc50 (wc50, n_125);
  or g631 (n_170, A[5], n_159, wc51);
  not gc51 (wc51, n_355);
  or g632 (n_386, n_320, wc52);
  not gc52 (wc52, n_177);
  or g633 (n_399, A[12], wc53);
  not gc53 (wc53, n_184);
  or g634 (n_196, A[9], wc54, wc55);
  not gc55 (wc55, n_176);
  not gc54 (wc54, n_406);
  xnor g635 (n_416, n_194, n_169);
  or g636 (n_417, n_169, wc56);
  not gc56 (wc56, n_194);
  xnor g637 (n_23, n_199, n_198);
  or g640 (n_455, wc57, n_208);
  not gc57 (wc57, n_68);
  xnor g641 (n_458, n_208, n_68);
  xnor g642 (n_180, n_384, n_320);
  or g643 (n_418, wc58, n_169);
  not gc58 (wc58, n_196);
  or g644 (n_50, n_198, wc59, n_199);
  not gc59 (wc59, n_422);
  or g645 (n_441, wc60, n_435);
  not gc60 (wc60, A[2]);
  or g646 (n_442, wc61, n_435);
  not gc61 (wc61, A[1]);
  xnor g647 (Z[2], n_435, n_443);
  or g648 (n_550, A[13], wc62);
  not gc62 (wc62, n_49);
  xnor g649 (n_553, n_49, A[13]);
  or g650 (n_456, wc63, n_208);
  not gc63 (wc63, n_454);
  or g651 (n_551, A[13], wc64);
  not gc64 (wc64, n_549);
  or g652 (n_557, A[14], wc65);
  not gc65 (wc65, n_554);
  xnor g653 (Z[25], n_316, n_554);
  or g654 (n_562, A[15], wc66);
  not gc66 (wc66, n_559);
  xnor g655 (Z[26], n_332, n_559);
endmodule

module mult_signed_const_751_GENERIC(A, Z);
  input [16:0] A;
  output [27:0] Z;
  wire [16:0] A;
  wire [27:0] Z;
  mult_signed_const_751_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

